LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE work.PIC_pkg.all;

entity ROM_Generated is
  port (
    Instruction     : out std_logic_vector(11 downto 0);
    Program_counter : in  std_logic_vector(11 downto 0));
end ROM_Generated;

architecture AUTOMATIC of ROM_Generated is
begin
    with Program_counter select
        Instruction <=
            X"0" & TYPE_2 & JMP_UNCOND when X"000",
            X"881" when X"001",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"002",
            X"000" when X"003",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"004",
            X"049" when X"005",
            X"0" & TYPE_1 & ALU_CMPE when X"006",
            X"0" & TYPE_2 & JMP_COND when X"007",
            X"00B" when X"008",
            X"0" & TYPE_2 & JMP_UNCOND when X"009",
            X"053" when X"00A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"00B",
            X"001" when X"00C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"00D",
            X"030" when X"00E",
            X"0" & TYPE_1 & ALU_SUB when X"00F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"010",
            X"043" when X"011",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"012",
            X"002" when X"013",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"014",
            X"030" when X"015",
            X"0" & TYPE_1 & ALU_SUB when X"016",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"017",
            X"044" when X"018",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"019",
            X"043" when X"01A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"01B",
            X"007" when X"01C",
            X"0" & TYPE_1 & ALU_CMPG when X"01D",
            X"0" & TYPE_2 & JMP_COND when X"01E",
            X"022" when X"01F",
            X"0" & TYPE_2 & JMP_UNCOND when X"020",
            X"02D" when X"021",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"022",
            X"045" when X"023",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"024",
            X"004" when X"025",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"026",
            X"052" when X"027",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"028",
            X"005" when X"029",
            X"0" & TYPE_4 & I_SEND when X"02A",
            X"0" & TYPE_2 & JMP_UNCOND when X"02B",
            X"880" when X"02C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"02D",
            X"044" when X"02E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"02F",
            X"001" when X"030",
            X"0" & TYPE_1 & ALU_CMPG when X"031",
            X"0" & TYPE_2 & JMP_COND when X"032",
            X"036" when X"033",
            X"0" & TYPE_2 & JMP_UNCOND when X"034",
            X"041" when X"035",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"036",
            X"045" when X"037",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"038",
            X"004" when X"039",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"03A",
            X"052" when X"03B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"03C",
            X"005" when X"03D",
            X"0" & TYPE_4 & I_SEND when X"03E",
            X"0" & TYPE_2 & JMP_UNCOND when X"03F",
            X"880" when X"040",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"041",
            X"043" when X"042",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"043",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"044",
            X"044" when X"045",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"046",
            X"010" when X"047",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"048",
            X"04F" when X"049",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"04A",
            X"004" when X"04B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"04C",
            X"04B" when X"04D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"04E",
            X"005" when X"04F",
            X"0" & TYPE_4 & I_SEND when X"050",
            X"0" & TYPE_2 & JMP_UNCOND when X"051",
            X"880" when X"052",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"053",
            X"000" when X"054",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"055",
            X"041" when X"056",
            X"0" & TYPE_1 & ALU_CMPE when X"057",
            X"0" & TYPE_2 & JMP_COND when X"058",
            X"05C" when X"059",
            X"0" & TYPE_2 & JMP_UNCOND when X"05A",
            X"0A4" when X"05B",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"05C",
            X"001" when X"05D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"05E",
            X"030" when X"05F",
            X"0" & TYPE_1 & ALU_SUB when X"060",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"061",
            X"043" when X"062",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"063",
            X"002" when X"064",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"065",
            X"030" when X"066",
            X"0" & TYPE_1 & ALU_SUB when X"067",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"068",
            X"044" when X"069",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"06A",
            X"043" when X"06B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"06C",
            X"009" when X"06D",
            X"0" & TYPE_1 & ALU_CMPG when X"06E",
            X"0" & TYPE_2 & JMP_COND when X"06F",
            X"073" when X"070",
            X"0" & TYPE_2 & JMP_UNCOND when X"071",
            X"07E" when X"072",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"073",
            X"045" when X"074",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"075",
            X"004" when X"076",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"077",
            X"052" when X"078",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"079",
            X"005" when X"07A",
            X"0" & TYPE_4 & I_SEND when X"07B",
            X"0" & TYPE_2 & JMP_UNCOND when X"07C",
            X"880" when X"07D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"07E",
            X"044" when X"07F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"080",
            X"009" when X"081",
            X"0" & TYPE_1 & ALU_CMPG when X"082",
            X"0" & TYPE_2 & JMP_COND when X"083",
            X"087" when X"084",
            X"0" & TYPE_2 & JMP_UNCOND when X"085",
            X"092" when X"086",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"087",
            X"045" when X"088",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"089",
            X"004" when X"08A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"08B",
            X"052" when X"08C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"08D",
            X"005" when X"08E",
            X"0" & TYPE_4 & I_SEND when X"08F",
            X"0" & TYPE_2 & JMP_UNCOND when X"090",
            X"880" when X"091",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"092",
            X"043" when X"093",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"094",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"095",
            X"044" when X"096",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"097",
            X"020" when X"098",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"099",
            X"04F" when X"09A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"09B",
            X"004" when X"09C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"09D",
            X"04B" when X"09E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"09F",
            X"005" when X"0A0",
            X"0" & TYPE_4 & I_SEND when X"0A1",
            X"0" & TYPE_2 & JMP_UNCOND when X"0A2",
            X"880" when X"0A3",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0A4",
            X"000" when X"0A5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0A6",
            X"054" when X"0A7",
            X"0" & TYPE_1 & ALU_CMPE when X"0A8",
            X"0" & TYPE_2 & JMP_COND when X"0A9",
            X"0AD" when X"0AA",
            X"0" & TYPE_2 & JMP_UNCOND when X"0AB",
            X"114" when X"0AC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0AD",
            X"001" when X"0AE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0AF",
            X"030" when X"0B0",
            X"0" & TYPE_1 & ALU_CMPL when X"0B1",
            X"0" & TYPE_2 & JMP_COND when X"0B2",
            X"0B6" when X"0B3",
            X"0" & TYPE_2 & JMP_UNCOND when X"0B4",
            X"0C1" when X"0B5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0B6",
            X"045" when X"0B7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0B8",
            X"004" when X"0B9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0BA",
            X"052" when X"0BB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0BC",
            X"005" when X"0BD",
            X"0" & TYPE_4 & I_SEND when X"0BE",
            X"0" & TYPE_2 & JMP_UNCOND when X"0BF",
            X"880" when X"0C0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0C1",
            X"001" when X"0C2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0C3",
            X"032" when X"0C4",
            X"0" & TYPE_1 & ALU_CMPG when X"0C5",
            X"0" & TYPE_2 & JMP_COND when X"0C6",
            X"0CA" when X"0C7",
            X"0" & TYPE_2 & JMP_UNCOND when X"0C8",
            X"0D5" when X"0C9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0CA",
            X"045" when X"0CB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0CC",
            X"004" when X"0CD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0CE",
            X"052" when X"0CF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0D0",
            X"005" when X"0D1",
            X"0" & TYPE_4 & I_SEND when X"0D2",
            X"0" & TYPE_2 & JMP_UNCOND when X"0D3",
            X"880" when X"0D4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0D5",
            X"002" when X"0D6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0D7",
            X"039" when X"0D8",
            X"0" & TYPE_1 & ALU_CMPG when X"0D9",
            X"0" & TYPE_2 & JMP_COND when X"0DA",
            X"0DE" when X"0DB",
            X"0" & TYPE_2 & JMP_UNCOND when X"0DC",
            X"0E9" when X"0DD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0DE",
            X"045" when X"0DF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0E0",
            X"004" when X"0E1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0E2",
            X"052" when X"0E3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0E4",
            X"005" when X"0E5",
            X"0" & TYPE_4 & I_SEND when X"0E6",
            X"0" & TYPE_2 & JMP_UNCOND when X"0E7",
            X"880" when X"0E8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0E9",
            X"001" when X"0EA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0EB",
            X"030" when X"0EC",
            X"0" & TYPE_1 & ALU_SUB when X"0ED",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0EE",
            X"045" when X"0EF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0F0",
            X"045" when X"0F1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0F2",
            X"000" when X"0F3",
            X"0" & TYPE_1 & ALU_ADD when X"0F4",
            X"0" & TYPE_1 & ALU_SHIFTL when X"0F5",
            X"0" & TYPE_1 & ALU_SHIFTL when X"0F6",
            X"0" & TYPE_1 & ALU_SHIFTL when X"0F7",
            X"0" & TYPE_1 & ALU_SHIFTL when X"0F8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0F9",
            X"045" when X"0FA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"0FB",
            X"002" when X"0FC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"0FD",
            X"030" when X"0FE",
            X"0" & TYPE_1 & ALU_SUB when X"0FF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"100",
            X"046" when X"101",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"102",
            X"045" when X"103",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"104",
            X"046" when X"105",
            X"0" & TYPE_1 & ALU_ADD when X"106",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"107",
            X"031" when X"108",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"109",
            X"04F" when X"10A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"10B",
            X"004" when X"10C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"10D",
            X"04B" when X"10E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"10F",
            X"005" when X"110",
            X"0" & TYPE_4 & I_SEND when X"111",
            X"0" & TYPE_2 & JMP_UNCOND when X"112",
            X"880" when X"113",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"114",
            X"000" when X"115",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"116",
            X"053" when X"117",
            X"0" & TYPE_1 & ALU_CMPE when X"118",
            X"0" & TYPE_2 & JMP_COND when X"119",
            X"11D" when X"11A",
            X"0" & TYPE_2 & JMP_UNCOND when X"11B",
            X"4A6" when X"11C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"11D",
            X"001" when X"11E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"11F",
            X"054" when X"120",
            X"0" & TYPE_1 & ALU_CMPE when X"121",
            X"0" & TYPE_2 & JMP_COND when X"122",
            X"126" when X"123",
            X"0" & TYPE_2 & JMP_UNCOND when X"124",
            X"147" when X"125",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"126",
            X"031" when X"127",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"128",
            X"000" when X"129",
            X"0" & TYPE_1 & ALU_ADD when X"12A",
            X"0" & TYPE_1 & ALU_SHIFTR when X"12B",
            X"0" & TYPE_1 & ALU_SHIFTR when X"12C",
            X"0" & TYPE_1 & ALU_SHIFTR when X"12D",
            X"0" & TYPE_1 & ALU_SHIFTR when X"12E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"12F",
            X"045" when X"130",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"131",
            X"031" when X"132",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"133",
            X"00F" when X"134",
            X"0" & TYPE_1 & ALU_AND when X"135",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"136",
            X"046" when X"137",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"138",
            X"045" when X"139",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"13A",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"13B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"13C",
            X"004" when X"13D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"13E",
            X"046" when X"13F",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"140",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"141",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"142",
            X"005" when X"143",
            X"0" & TYPE_4 & I_SEND when X"144",
            X"0" & TYPE_2 & JMP_UNCOND when X"145",
            X"880" when X"146",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"147",
            X"001" when X"148",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"149",
            X"041" when X"14A",
            X"0" & TYPE_1 & ALU_CMPE when X"14B",
            X"0" & TYPE_2 & JMP_COND when X"14C",
            X"150" when X"14D",
            X"0" & TYPE_2 & JMP_UNCOND when X"14E",
            X"17F" when X"14F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"150",
            X"002" when X"151",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"152",
            X"030" when X"153",
            X"0" & TYPE_1 & ALU_SUB when X"154",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"155",
            X"043" when X"156",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"157",
            X"043" when X"158",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"159",
            X"009" when X"15A",
            X"0" & TYPE_1 & ALU_CMPG when X"15B",
            X"0" & TYPE_2 & JMP_COND when X"15C",
            X"160" when X"15D",
            X"0" & TYPE_2 & JMP_UNCOND when X"15E",
            X"16B" when X"15F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"160",
            X"045" when X"161",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"162",
            X"004" when X"163",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"164",
            X"052" when X"165",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"166",
            X"005" when X"167",
            X"0" & TYPE_4 & I_SEND when X"168",
            X"0" & TYPE_2 & JMP_UNCOND when X"169",
            X"880" when X"16A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"16B",
            X"043" when X"16C",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"16D",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"16E",
            X"020" when X"16F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"170",
            X"044" when X"171",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"172",
            X"041" when X"173",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"174",
            X"004" when X"175",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"176",
            X"044" when X"177",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"178",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"179",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"17A",
            X"005" when X"17B",
            X"0" & TYPE_4 & I_SEND when X"17C",
            X"0" & TYPE_2 & JMP_UNCOND when X"17D",
            X"880" when X"17E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"17F",
            X"001" when X"180",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"181",
            X"049" when X"182",
            X"0" & TYPE_1 & ALU_CMPE when X"183",
            X"0" & TYPE_2 & JMP_COND when X"184",
            X"188" when X"185",
            X"0" & TYPE_2 & JMP_UNCOND when X"186",
            X"1B7" when X"187",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"188",
            X"002" when X"189",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"18A",
            X"030" when X"18B",
            X"0" & TYPE_1 & ALU_SUB when X"18C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"18D",
            X"043" when X"18E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"18F",
            X"043" when X"190",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"191",
            X"007" when X"192",
            X"0" & TYPE_1 & ALU_CMPG when X"193",
            X"0" & TYPE_2 & JMP_COND when X"194",
            X"198" when X"195",
            X"0" & TYPE_2 & JMP_UNCOND when X"196",
            X"1A3" when X"197",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"198",
            X"045" when X"199",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"19A",
            X"004" when X"19B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"19C",
            X"052" when X"19D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"19E",
            X"005" when X"19F",
            X"0" & TYPE_4 & I_SEND when X"1A0",
            X"0" & TYPE_2 & JMP_UNCOND when X"1A1",
            X"880" when X"1A2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1A3",
            X"043" when X"1A4",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"1A5",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"1A6",
            X"010" when X"1A7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1A8",
            X"044" when X"1A9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1AA",
            X"049" when X"1AB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1AC",
            X"004" when X"1AD",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1AE",
            X"044" when X"1AF",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"1B0",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"1B1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1B2",
            X"005" when X"1B3",
            X"0" & TYPE_4 & I_SEND when X"1B4",
            X"0" & TYPE_2 & JMP_UNCOND when X"1B5",
            X"880" when X"1B6",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1B7",
            X"001" when X"1B8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"1B9",
            X"052" when X"1BA",
            X"0" & TYPE_1 & ALU_CMPE when X"1BB",
            X"0" & TYPE_2 & JMP_COND when X"1BC",
            X"1C0" when X"1BD",
            X"0" & TYPE_2 & JMP_UNCOND when X"1BE",
            X"4A6" when X"1BF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1C0",
            X"042" when X"1C1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1C2",
            X"004" when X"1C3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1C4",
            X"041" when X"1C5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1C6",
            X"005" when X"1C7",
            X"0" & TYPE_4 & I_SEND when X"1C8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1C9",
            X"055" when X"1CA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1CB",
            X"004" when X"1CC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1CD",
            X"044" when X"1CE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1CF",
            X"005" when X"1D0",
            X"0" & TYPE_4 & I_SEND when X"1D1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1D2",
            X"03A" when X"1D3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1D4",
            X"004" when X"1D5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1D6",
            X"020" when X"1D7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1D8",
            X"005" when X"1D9",
            X"0" & TYPE_4 & I_SEND when X"1DA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1DB",
            X"009" when X"1DC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"1DD",
            X"000" when X"1DE",
            X"0" & TYPE_1 & ALU_CMPE when X"1DF",
            X"0" & TYPE_2 & JMP_COND when X"1E0",
            X"1E4" when X"1E1",
            X"0" & TYPE_2 & JMP_UNCOND when X"1E2",
            X"1F6" when X"1E3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1E4",
            X"033" when X"1E5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1E6",
            X"004" when X"1E7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1E8",
            X"030" when X"1E9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1EA",
            X"005" when X"1EB",
            X"0" & TYPE_4 & I_SEND when X"1EC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1ED",
            X"030" when X"1EE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1EF",
            X"004" when X"1F0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1F1",
            X"020" when X"1F2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1F3",
            X"005" when X"1F4",
            X"0" & TYPE_4 & I_SEND when X"1F5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1F6",
            X"009" when X"1F7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"1F8",
            X"001" when X"1F9",
            X"0" & TYPE_1 & ALU_CMPE when X"1FA",
            X"0" & TYPE_2 & JMP_COND when X"1FB",
            X"1FF" when X"1FC",
            X"0" & TYPE_2 & JMP_UNCOND when X"1FD",
            X"21A" when X"1FE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1FF",
            X"031" when X"200",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"201",
            X"004" when X"202",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"203",
            X"032" when X"204",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"205",
            X"005" when X"206",
            X"0" & TYPE_4 & I_SEND when X"207",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"208",
            X"030" when X"209",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"20A",
            X"004" when X"20B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"20C",
            X"030" when X"20D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"20E",
            X"005" when X"20F",
            X"0" & TYPE_4 & I_SEND when X"210",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"211",
            X"020" when X"212",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"213",
            X"004" when X"214",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"215",
            X"020" when X"216",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"217",
            X"005" when X"218",
            X"0" & TYPE_4 & I_SEND when X"219",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"21A",
            X"009" when X"21B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"21C",
            X"002" when X"21D",
            X"0" & TYPE_1 & ALU_CMPE when X"21E",
            X"0" & TYPE_2 & JMP_COND when X"21F",
            X"223" when X"220",
            X"0" & TYPE_2 & JMP_UNCOND when X"221",
            X"23E" when X"222",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"223",
            X"032" when X"224",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"225",
            X"004" when X"226",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"227",
            X"034" when X"228",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"229",
            X"005" when X"22A",
            X"0" & TYPE_4 & I_SEND when X"22B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"22C",
            X"030" when X"22D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"22E",
            X"004" when X"22F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"230",
            X"030" when X"231",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"232",
            X"005" when X"233",
            X"0" & TYPE_4 & I_SEND when X"234",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"235",
            X"020" when X"236",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"237",
            X"004" when X"238",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"239",
            X"020" when X"23A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"23B",
            X"005" when X"23C",
            X"0" & TYPE_4 & I_SEND when X"23D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"23E",
            X"009" when X"23F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"240",
            X"003" when X"241",
            X"0" & TYPE_1 & ALU_CMPE when X"242",
            X"0" & TYPE_2 & JMP_COND when X"243",
            X"247" when X"244",
            X"0" & TYPE_2 & JMP_UNCOND when X"245",
            X"262" when X"246",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"247",
            X"034" when X"248",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"249",
            X"004" when X"24A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"24B",
            X"038" when X"24C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"24D",
            X"005" when X"24E",
            X"0" & TYPE_4 & I_SEND when X"24F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"250",
            X"030" when X"251",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"252",
            X"004" when X"253",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"254",
            X"030" when X"255",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"256",
            X"005" when X"257",
            X"0" & TYPE_4 & I_SEND when X"258",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"259",
            X"020" when X"25A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"25B",
            X"004" when X"25C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"25D",
            X"020" when X"25E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"25F",
            X"005" when X"260",
            X"0" & TYPE_4 & I_SEND when X"261",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"262",
            X"009" when X"263",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"264",
            X"004" when X"265",
            X"0" & TYPE_1 & ALU_CMPE when X"266",
            X"0" & TYPE_2 & JMP_COND when X"267",
            X"26B" when X"268",
            X"0" & TYPE_2 & JMP_UNCOND when X"269",
            X"286" when X"26A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"26B",
            X"039" when X"26C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"26D",
            X"004" when X"26E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"26F",
            X"036" when X"270",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"271",
            X"005" when X"272",
            X"0" & TYPE_4 & I_SEND when X"273",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"274",
            X"030" when X"275",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"276",
            X"004" when X"277",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"278",
            X"030" when X"279",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"27A",
            X"005" when X"27B",
            X"0" & TYPE_4 & I_SEND when X"27C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"27D",
            X"020" when X"27E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"27F",
            X"004" when X"280",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"281",
            X"020" when X"282",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"283",
            X"005" when X"284",
            X"0" & TYPE_4 & I_SEND when X"285",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"286",
            X"009" when X"287",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"288",
            X"005" when X"289",
            X"0" & TYPE_1 & ALU_CMPE when X"28A",
            X"0" & TYPE_2 & JMP_COND when X"28B",
            X"28F" when X"28C",
            X"0" & TYPE_2 & JMP_UNCOND when X"28D",
            X"2AA" when X"28E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"28F",
            X"031" when X"290",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"291",
            X"004" when X"292",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"293",
            X"039" when X"294",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"295",
            X"005" when X"296",
            X"0" & TYPE_4 & I_SEND when X"297",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"298",
            X"032" when X"299",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"29A",
            X"004" when X"29B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"29C",
            X"030" when X"29D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"29E",
            X"005" when X"29F",
            X"0" & TYPE_4 & I_SEND when X"2A0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2A1",
            X"030" when X"2A2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2A3",
            X"004" when X"2A4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2A5",
            X"020" when X"2A6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2A7",
            X"005" when X"2A8",
            X"0" & TYPE_4 & I_SEND when X"2A9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"2AA",
            X"009" when X"2AB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"2AC",
            X"006" when X"2AD",
            X"0" & TYPE_1 & ALU_CMPE when X"2AE",
            X"0" & TYPE_2 & JMP_COND when X"2AF",
            X"2B3" when X"2B0",
            X"0" & TYPE_2 & JMP_UNCOND when X"2B1",
            X"2CE" when X"2B2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2B3",
            X"033" when X"2B4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2B5",
            X"004" when X"2B6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2B7",
            X"038" when X"2B8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2B9",
            X"005" when X"2BA",
            X"0" & TYPE_4 & I_SEND when X"2BB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2BC",
            X"034" when X"2BD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2BE",
            X"004" when X"2BF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2C0",
            X"030" when X"2C1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2C2",
            X"005" when X"2C3",
            X"0" & TYPE_4 & I_SEND when X"2C4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2C5",
            X"030" when X"2C6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2C7",
            X"004" when X"2C8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2C9",
            X"020" when X"2CA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2CB",
            X"005" when X"2CC",
            X"0" & TYPE_4 & I_SEND when X"2CD",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"2CE",
            X"009" when X"2CF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"2D0",
            X"007" when X"2D1",
            X"0" & TYPE_1 & ALU_CMPE when X"2D2",
            X"0" & TYPE_2 & JMP_COND when X"2D3",
            X"2D7" when X"2D4",
            X"0" & TYPE_2 & JMP_UNCOND when X"2D5",
            X"2F2" when X"2D6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2D7",
            X"035" when X"2D8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2D9",
            X"004" when X"2DA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2DB",
            X"037" when X"2DC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2DD",
            X"005" when X"2DE",
            X"0" & TYPE_4 & I_SEND when X"2DF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2E0",
            X"036" when X"2E1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2E2",
            X"004" when X"2E3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2E4",
            X"030" when X"2E5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2E6",
            X"005" when X"2E7",
            X"0" & TYPE_4 & I_SEND when X"2E8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2E9",
            X"030" when X"2EA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2EB",
            X"004" when X"2EC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2ED",
            X"020" when X"2EE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2EF",
            X"005" when X"2F0",
            X"0" & TYPE_4 & I_SEND when X"2F1",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"2F2",
            X"009" when X"2F3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"2F4",
            X"008" when X"2F5",
            X"0" & TYPE_1 & ALU_CMPE when X"2F6",
            X"0" & TYPE_2 & JMP_COND when X"2F7",
            X"2FB" when X"2F8",
            X"0" & TYPE_2 & JMP_UNCOND when X"2F9",
            X"31F" when X"2FA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2FB",
            X"031" when X"2FC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"2FD",
            X"004" when X"2FE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"2FF",
            X"031" when X"300",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"301",
            X"005" when X"302",
            X"0" & TYPE_4 & I_SEND when X"303",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"304",
            X"035" when X"305",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"306",
            X"004" when X"307",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"308",
            X"032" when X"309",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"30A",
            X"005" when X"30B",
            X"0" & TYPE_4 & I_SEND when X"30C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"30D",
            X"030" when X"30E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"30F",
            X"004" when X"310",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"311",
            X"030" when X"312",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"313",
            X"005" when X"314",
            X"0" & TYPE_4 & I_SEND when X"315",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"316",
            X"020" when X"317",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"318",
            X"004" when X"319",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"31A",
            X"020" when X"31B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"31C",
            X"005" when X"31D",
            X"0" & TYPE_4 & I_SEND when X"31E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"31F",
            X"009" when X"320",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"321",
            X"009" when X"322",
            X"0" & TYPE_1 & ALU_CMPE when X"323",
            X"0" & TYPE_2 & JMP_COND when X"324",
            X"328" when X"325",
            X"0" & TYPE_2 & JMP_UNCOND when X"326",
            X"34C" when X"327",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"328",
            X"032" when X"329",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"32A",
            X"004" when X"32B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"32C",
            X"033" when X"32D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"32E",
            X"005" when X"32F",
            X"0" & TYPE_4 & I_SEND when X"330",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"331",
            X"030" when X"332",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"333",
            X"004" when X"334",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"335",
            X"034" when X"336",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"337",
            X"005" when X"338",
            X"0" & TYPE_4 & I_SEND when X"339",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"33A",
            X"030" when X"33B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"33C",
            X"004" when X"33D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"33E",
            X"030" when X"33F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"340",
            X"005" when X"341",
            X"0" & TYPE_4 & I_SEND when X"342",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"343",
            X"020" when X"344",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"345",
            X"004" when X"346",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"347",
            X"020" when X"348",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"349",
            X"005" when X"34A",
            X"0" & TYPE_4 & I_SEND when X"34B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"34C",
            X"04E" when X"34D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"34E",
            X"004" when X"34F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"350",
            X"05F" when X"351",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"352",
            X"005" when X"353",
            X"0" & TYPE_4 & I_SEND when X"354",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"355",
            X"042" when X"356",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"357",
            X"004" when X"358",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"359",
            X"049" when X"35A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"35B",
            X"005" when X"35C",
            X"0" & TYPE_4 & I_SEND when X"35D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"35E",
            X"054" when X"35F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"360",
            X"004" when X"361",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"362",
            X"053" when X"363",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"364",
            X"005" when X"365",
            X"0" & TYPE_4 & I_SEND when X"366",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"367",
            X"03A" when X"368",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"369",
            X"004" when X"36A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"36B",
            X"020" when X"36C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"36D",
            X"005" when X"36E",
            X"0" & TYPE_4 & I_SEND when X"36F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"370",
            X"008" when X"371",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"372",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"373",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"374",
            X"004" when X"375",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"376",
            X"020" when X"377",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"378",
            X"005" when X"379",
            X"0" & TYPE_4 & I_SEND when X"37A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"37B",
            X"053" when X"37C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"37D",
            X"004" when X"37E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"37F",
            X"054" when X"380",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"381",
            X"005" when X"382",
            X"0" & TYPE_4 & I_SEND when X"383",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"384",
            X"04F" when X"385",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"386",
            X"004" when X"387",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"388",
            X"050" when X"389",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"38A",
            X"005" when X"38B",
            X"0" & TYPE_4 & I_SEND when X"38C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"38D",
            X"03A" when X"38E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"38F",
            X"004" when X"390",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"391",
            X"020" when X"392",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"393",
            X"005" when X"394",
            X"0" & TYPE_4 & I_SEND when X"395",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"396",
            X"007" when X"397",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"398",
            X"002" when X"399",
            X"0" & TYPE_1 & ALU_CMPE when X"39A",
            X"0" & TYPE_2 & JMP_COND when X"39B",
            X"39F" when X"39C",
            X"0" & TYPE_2 & JMP_UNCOND when X"39D",
            X"3A8" when X"39E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"39F",
            X"031" when X"3A0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3A1",
            X"004" when X"3A2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3A3",
            X"020" when X"3A4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3A5",
            X"005" when X"3A6",
            X"0" & TYPE_4 & I_SEND when X"3A7",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"3A8",
            X"007" when X"3A9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"3AA",
            X"003" when X"3AB",
            X"0" & TYPE_1 & ALU_CMPE when X"3AC",
            X"0" & TYPE_2 & JMP_COND when X"3AD",
            X"3B1" when X"3AE",
            X"0" & TYPE_2 & JMP_UNCOND when X"3AF",
            X"3C3" when X"3B0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3B1",
            X"031" when X"3B2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3B3",
            X"004" when X"3B4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3B5",
            X"02E" when X"3B6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3B7",
            X"005" when X"3B8",
            X"0" & TYPE_4 & I_SEND when X"3B9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3BA",
            X"035" when X"3BB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3BC",
            X"004" when X"3BD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3BE",
            X"020" when X"3BF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3C0",
            X"005" when X"3C1",
            X"0" & TYPE_4 & I_SEND when X"3C2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"3C3",
            X"007" when X"3C4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"3C5",
            X"004" when X"3C6",
            X"0" & TYPE_1 & ALU_CMPE when X"3C7",
            X"0" & TYPE_2 & JMP_COND when X"3C8",
            X"3CC" when X"3C9",
            X"0" & TYPE_2 & JMP_UNCOND when X"3CA",
            X"3D5" when X"3CB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3CC",
            X"032" when X"3CD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3CE",
            X"004" when X"3CF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3D0",
            X"020" when X"3D1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3D2",
            X"005" when X"3D3",
            X"0" & TYPE_4 & I_SEND when X"3D4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3D5",
            X"050" when X"3D6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3D7",
            X"004" when X"3D8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3D9",
            X"041" when X"3DA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3DB",
            X"005" when X"3DC",
            X"0" & TYPE_4 & I_SEND when X"3DD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3DE",
            X"052" when X"3DF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3E0",
            X"004" when X"3E1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3E2",
            X"049" when X"3E3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3E4",
            X"005" when X"3E5",
            X"0" & TYPE_4 & I_SEND when X"3E6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3E7",
            X"054" when X"3E8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3E9",
            X"004" when X"3EA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3EB",
            X"059" when X"3EC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3ED",
            X"005" when X"3EE",
            X"0" & TYPE_4 & I_SEND when X"3EF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3F0",
            X"03A" when X"3F1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3F2",
            X"004" when X"3F3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"3F4",
            X"020" when X"3F5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"3F6",
            X"005" when X"3F7",
            X"0" & TYPE_4 & I_SEND when X"3F8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"3F9",
            X"050" when X"3FA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"3FB",
            X"000" when X"3FC",
            X"0" & TYPE_1 & ALU_CMPE when X"3FD",
            X"0" & TYPE_2 & JMP_COND when X"3FE",
            X"402" when X"3FF",
            X"0" & TYPE_2 & JMP_UNCOND when X"400",
            X"41D" when X"401",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"402",
            X"045" when X"403",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"404",
            X"004" when X"405",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"406",
            X"056" when X"407",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"408",
            X"005" when X"409",
            X"0" & TYPE_4 & I_SEND when X"40A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"40B",
            X"045" when X"40C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"40D",
            X"004" when X"40E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"40F",
            X"04E" when X"410",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"411",
            X"005" when X"412",
            X"0" & TYPE_4 & I_SEND when X"413",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"414",
            X"020" when X"415",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"416",
            X"004" when X"417",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"418",
            X"020" when X"419",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"41A",
            X"005" when X"41B",
            X"0" & TYPE_4 & I_SEND when X"41C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"41D",
            X"050" when X"41E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"41F",
            X"001" when X"420",
            X"0" & TYPE_1 & ALU_CMPE when X"421",
            X"0" & TYPE_2 & JMP_COND when X"422",
            X"426" when X"423",
            X"0" & TYPE_2 & JMP_UNCOND when X"424",
            X"438" when X"425",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"426",
            X"04F" when X"427",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"428",
            X"004" when X"429",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"42A",
            X"044" when X"42B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"42C",
            X"005" when X"42D",
            X"0" & TYPE_4 & I_SEND when X"42E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"42F",
            X"044" when X"430",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"431",
            X"004" when X"432",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"433",
            X"020" when X"434",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"435",
            X"005" when X"436",
            X"0" & TYPE_4 & I_SEND when X"437",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"438",
            X"050" when X"439",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"43A",
            X"002" when X"43B",
            X"0" & TYPE_1 & ALU_CMPE when X"43C",
            X"0" & TYPE_2 & JMP_COND when X"43D",
            X"441" when X"43E",
            X"0" & TYPE_2 & JMP_UNCOND when X"43F",
            X"45C" when X"440",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"441",
            X"04D" when X"442",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"443",
            X"004" when X"444",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"445",
            X"041" when X"446",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"447",
            X"005" when X"448",
            X"0" & TYPE_4 & I_SEND when X"449",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"44A",
            X"052" when X"44B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"44C",
            X"004" when X"44D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"44E",
            X"04B" when X"44F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"450",
            X"005" when X"451",
            X"0" & TYPE_4 & I_SEND when X"452",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"453",
            X"020" when X"454",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"455",
            X"004" when X"456",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"457",
            X"020" when X"458",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"459",
            X"005" when X"45A",
            X"0" & TYPE_4 & I_SEND when X"45B",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"45C",
            X"050" when X"45D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"45E",
            X"003" when X"45F",
            X"0" & TYPE_1 & ALU_CMPE when X"460",
            X"0" & TYPE_2 & JMP_COND when X"461",
            X"465" when X"462",
            X"0" & TYPE_2 & JMP_UNCOND when X"463",
            X"480" when X"464",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"465",
            X"053" when X"466",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"467",
            X"004" when X"468",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"469",
            X"050" when X"46A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"46B",
            X"005" when X"46C",
            X"0" & TYPE_4 & I_SEND when X"46D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"46E",
            X"041" when X"46F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"470",
            X"004" when X"471",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"472",
            X"043" when X"473",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"474",
            X"005" when X"475",
            X"0" & TYPE_4 & I_SEND when X"476",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"477",
            X"045" when X"478",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"479",
            X"004" when X"47A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"47B",
            X"020" when X"47C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"47D",
            X"005" when X"47E",
            X"0" & TYPE_4 & I_SEND when X"47F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"480",
            X"050" when X"481",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"482",
            X"004" when X"483",
            X"0" & TYPE_1 & ALU_CMPE when X"484",
            X"0" & TYPE_2 & JMP_COND when X"485",
            X"489" when X"486",
            X"0" & TYPE_2 & JMP_UNCOND when X"487",
            X"4A4" when X"488",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"489",
            X"04E" when X"48A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"48B",
            X"004" when X"48C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"48D",
            X"04F" when X"48E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"48F",
            X"005" when X"490",
            X"0" & TYPE_4 & I_SEND when X"491",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"492",
            X"04E" when X"493",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"494",
            X"004" when X"495",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"496",
            X"045" when X"497",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"498",
            X"005" when X"499",
            X"0" & TYPE_4 & I_SEND when X"49A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"49B",
            X"020" when X"49C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"49D",
            X"004" when X"49E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"49F",
            X"020" when X"4A0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4A1",
            X"005" when X"4A2",
            X"0" & TYPE_4 & I_SEND when X"4A3",
            X"0" & TYPE_2 & JMP_UNCOND when X"4A4",
            X"880" when X"4A5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"4A6",
            X"000" when X"4A7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"4A8",
            X"052" when X"4A9",
            X"0" & TYPE_1 & ALU_CMPE when X"4AA",
            X"0" & TYPE_2 & JMP_COND when X"4AB",
            X"4AF" when X"4AC",
            X"0" & TYPE_2 & JMP_UNCOND when X"4AD",
            X"880" when X"4AE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"4AF",
            X"002" when X"4B0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"4B1",
            X"030" when X"4B2",
            X"0" & TYPE_1 & ALU_SUB when X"4B3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4B4",
            X"044" when X"4B5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"4B6",
            X"001" when X"4B7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"4B8",
            X"039" when X"4B9",
            X"0" & TYPE_1 & ALU_CMPE when X"4BA",
            X"0" & TYPE_2 & JMP_COND when X"4BB",
            X"4BF" when X"4BC",
            X"0" & TYPE_2 & JMP_UNCOND when X"4BD",
            X"66E" when X"4BE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"4BF",
            X"044" when X"4C0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"4C1",
            X"009" when X"4C2",
            X"0" & TYPE_1 & ALU_CMPG when X"4C3",
            X"0" & TYPE_2 & JMP_COND when X"4C4",
            X"4C8" when X"4C5",
            X"0" & TYPE_2 & JMP_UNCOND when X"4C6",
            X"4D3" when X"4C7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4C8",
            X"045" when X"4C9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4CA",
            X"004" when X"4CB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4CC",
            X"052" when X"4CD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4CE",
            X"005" when X"4CF",
            X"0" & TYPE_4 & I_SEND when X"4D0",
            X"0" & TYPE_2 & JMP_UNCOND when X"4D1",
            X"880" when X"4D2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4D3",
            X"042" when X"4D4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4D5",
            X"004" when X"4D6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4D7",
            X"041" when X"4D8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4D9",
            X"005" when X"4DA",
            X"0" & TYPE_4 & I_SEND when X"4DB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4DC",
            X"055" when X"4DD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4DE",
            X"004" when X"4DF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4E0",
            X"044" when X"4E1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4E2",
            X"005" when X"4E3",
            X"0" & TYPE_4 & I_SEND when X"4E4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4E5",
            X"03A" when X"4E6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4E7",
            X"004" when X"4E8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4E9",
            X"020" when X"4EA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4EB",
            X"005" when X"4EC",
            X"0" & TYPE_4 & I_SEND when X"4ED",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"4EE",
            X"002" when X"4EF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"4F0",
            X"030" when X"4F1",
            X"0" & TYPE_1 & ALU_CMPE when X"4F2",
            X"0" & TYPE_2 & JMP_COND when X"4F3",
            X"4F7" when X"4F4",
            X"0" & TYPE_2 & JMP_UNCOND when X"4F5",
            X"509" when X"4F6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4F7",
            X"033" when X"4F8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4F9",
            X"004" when X"4FA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"4FB",
            X"030" when X"4FC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"4FD",
            X"005" when X"4FE",
            X"0" & TYPE_4 & I_SEND when X"4FF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"500",
            X"030" when X"501",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"502",
            X"004" when X"503",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"504",
            X"020" when X"505",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"506",
            X"005" when X"507",
            X"0" & TYPE_4 & I_SEND when X"508",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"509",
            X"002" when X"50A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"50B",
            X"031" when X"50C",
            X"0" & TYPE_1 & ALU_CMPE when X"50D",
            X"0" & TYPE_2 & JMP_COND when X"50E",
            X"512" when X"50F",
            X"0" & TYPE_2 & JMP_UNCOND when X"510",
            X"52D" when X"511",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"512",
            X"031" when X"513",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"514",
            X"004" when X"515",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"516",
            X"032" when X"517",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"518",
            X"005" when X"519",
            X"0" & TYPE_4 & I_SEND when X"51A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"51B",
            X"030" when X"51C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"51D",
            X"004" when X"51E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"51F",
            X"030" when X"520",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"521",
            X"005" when X"522",
            X"0" & TYPE_4 & I_SEND when X"523",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"524",
            X"020" when X"525",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"526",
            X"004" when X"527",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"528",
            X"020" when X"529",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"52A",
            X"005" when X"52B",
            X"0" & TYPE_4 & I_SEND when X"52C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"52D",
            X"002" when X"52E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"52F",
            X"032" when X"530",
            X"0" & TYPE_1 & ALU_CMPE when X"531",
            X"0" & TYPE_2 & JMP_COND when X"532",
            X"536" when X"533",
            X"0" & TYPE_2 & JMP_UNCOND when X"534",
            X"551" when X"535",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"536",
            X"032" when X"537",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"538",
            X"004" when X"539",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"53A",
            X"034" when X"53B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"53C",
            X"005" when X"53D",
            X"0" & TYPE_4 & I_SEND when X"53E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"53F",
            X"030" when X"540",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"541",
            X"004" when X"542",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"543",
            X"030" when X"544",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"545",
            X"005" when X"546",
            X"0" & TYPE_4 & I_SEND when X"547",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"548",
            X"020" when X"549",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"54A",
            X"004" when X"54B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"54C",
            X"020" when X"54D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"54E",
            X"005" when X"54F",
            X"0" & TYPE_4 & I_SEND when X"550",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"551",
            X"002" when X"552",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"553",
            X"033" when X"554",
            X"0" & TYPE_1 & ALU_CMPE when X"555",
            X"0" & TYPE_2 & JMP_COND when X"556",
            X"55A" when X"557",
            X"0" & TYPE_2 & JMP_UNCOND when X"558",
            X"575" when X"559",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"55A",
            X"034" when X"55B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"55C",
            X"004" when X"55D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"55E",
            X"038" when X"55F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"560",
            X"005" when X"561",
            X"0" & TYPE_4 & I_SEND when X"562",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"563",
            X"030" when X"564",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"565",
            X"004" when X"566",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"567",
            X"030" when X"568",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"569",
            X"005" when X"56A",
            X"0" & TYPE_4 & I_SEND when X"56B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"56C",
            X"020" when X"56D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"56E",
            X"004" when X"56F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"570",
            X"020" when X"571",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"572",
            X"005" when X"573",
            X"0" & TYPE_4 & I_SEND when X"574",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"575",
            X"002" when X"576",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"577",
            X"034" when X"578",
            X"0" & TYPE_1 & ALU_CMPE when X"579",
            X"0" & TYPE_2 & JMP_COND when X"57A",
            X"57E" when X"57B",
            X"0" & TYPE_2 & JMP_UNCOND when X"57C",
            X"599" when X"57D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"57E",
            X"039" when X"57F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"580",
            X"004" when X"581",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"582",
            X"036" when X"583",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"584",
            X"005" when X"585",
            X"0" & TYPE_4 & I_SEND when X"586",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"587",
            X"030" when X"588",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"589",
            X"004" when X"58A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"58B",
            X"030" when X"58C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"58D",
            X"005" when X"58E",
            X"0" & TYPE_4 & I_SEND when X"58F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"590",
            X"020" when X"591",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"592",
            X"004" when X"593",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"594",
            X"020" when X"595",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"596",
            X"005" when X"597",
            X"0" & TYPE_4 & I_SEND when X"598",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"599",
            X"002" when X"59A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"59B",
            X"035" when X"59C",
            X"0" & TYPE_1 & ALU_CMPE when X"59D",
            X"0" & TYPE_2 & JMP_COND when X"59E",
            X"5A2" when X"59F",
            X"0" & TYPE_2 & JMP_UNCOND when X"5A0",
            X"5BD" when X"5A1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5A2",
            X"031" when X"5A3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5A4",
            X"004" when X"5A5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5A6",
            X"039" when X"5A7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5A8",
            X"005" when X"5A9",
            X"0" & TYPE_4 & I_SEND when X"5AA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5AB",
            X"032" when X"5AC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5AD",
            X"004" when X"5AE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5AF",
            X"030" when X"5B0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5B1",
            X"005" when X"5B2",
            X"0" & TYPE_4 & I_SEND when X"5B3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5B4",
            X"030" when X"5B5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5B6",
            X"004" when X"5B7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5B8",
            X"020" when X"5B9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5BA",
            X"005" when X"5BB",
            X"0" & TYPE_4 & I_SEND when X"5BC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"5BD",
            X"002" when X"5BE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"5BF",
            X"036" when X"5C0",
            X"0" & TYPE_1 & ALU_CMPE when X"5C1",
            X"0" & TYPE_2 & JMP_COND when X"5C2",
            X"5C6" when X"5C3",
            X"0" & TYPE_2 & JMP_UNCOND when X"5C4",
            X"5E1" when X"5C5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5C6",
            X"033" when X"5C7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5C8",
            X"004" when X"5C9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5CA",
            X"038" when X"5CB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5CC",
            X"005" when X"5CD",
            X"0" & TYPE_4 & I_SEND when X"5CE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5CF",
            X"034" when X"5D0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5D1",
            X"004" when X"5D2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5D3",
            X"030" when X"5D4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5D5",
            X"005" when X"5D6",
            X"0" & TYPE_4 & I_SEND when X"5D7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5D8",
            X"030" when X"5D9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5DA",
            X"004" when X"5DB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5DC",
            X"020" when X"5DD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5DE",
            X"005" when X"5DF",
            X"0" & TYPE_4 & I_SEND when X"5E0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"5E1",
            X"002" when X"5E2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"5E3",
            X"037" when X"5E4",
            X"0" & TYPE_1 & ALU_CMPE when X"5E5",
            X"0" & TYPE_2 & JMP_COND when X"5E6",
            X"5EA" when X"5E7",
            X"0" & TYPE_2 & JMP_UNCOND when X"5E8",
            X"605" when X"5E9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5EA",
            X"035" when X"5EB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5EC",
            X"004" when X"5ED",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5EE",
            X"037" when X"5EF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5F0",
            X"005" when X"5F1",
            X"0" & TYPE_4 & I_SEND when X"5F2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5F3",
            X"036" when X"5F4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5F5",
            X"004" when X"5F6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5F7",
            X"030" when X"5F8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5F9",
            X"005" when X"5FA",
            X"0" & TYPE_4 & I_SEND when X"5FB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"5FC",
            X"030" when X"5FD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"5FE",
            X"004" when X"5FF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"600",
            X"020" when X"601",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"602",
            X"005" when X"603",
            X"0" & TYPE_4 & I_SEND when X"604",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"605",
            X"002" when X"606",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"607",
            X"038" when X"608",
            X"0" & TYPE_1 & ALU_CMPE when X"609",
            X"0" & TYPE_2 & JMP_COND when X"60A",
            X"60E" when X"60B",
            X"0" & TYPE_2 & JMP_UNCOND when X"60C",
            X"632" when X"60D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"60E",
            X"031" when X"60F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"610",
            X"004" when X"611",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"612",
            X"031" when X"613",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"614",
            X"005" when X"615",
            X"0" & TYPE_4 & I_SEND when X"616",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"617",
            X"035" when X"618",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"619",
            X"004" when X"61A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"61B",
            X"032" when X"61C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"61D",
            X"005" when X"61E",
            X"0" & TYPE_4 & I_SEND when X"61F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"620",
            X"030" when X"621",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"622",
            X"004" when X"623",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"624",
            X"030" when X"625",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"626",
            X"005" when X"627",
            X"0" & TYPE_4 & I_SEND when X"628",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"629",
            X"020" when X"62A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"62B",
            X"004" when X"62C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"62D",
            X"020" when X"62E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"62F",
            X"005" when X"630",
            X"0" & TYPE_4 & I_SEND when X"631",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"632",
            X"002" when X"633",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"634",
            X"039" when X"635",
            X"0" & TYPE_1 & ALU_CMPE when X"636",
            X"0" & TYPE_2 & JMP_COND when X"637",
            X"63B" when X"638",
            X"0" & TYPE_2 & JMP_UNCOND when X"639",
            X"65F" when X"63A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"63B",
            X"032" when X"63C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"63D",
            X"004" when X"63E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"63F",
            X"033" when X"640",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"641",
            X"005" when X"642",
            X"0" & TYPE_4 & I_SEND when X"643",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"644",
            X"030" when X"645",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"646",
            X"004" when X"647",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"648",
            X"034" when X"649",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"64A",
            X"005" when X"64B",
            X"0" & TYPE_4 & I_SEND when X"64C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"64D",
            X"030" when X"64E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"64F",
            X"004" when X"650",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"651",
            X"030" when X"652",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"653",
            X"005" when X"654",
            X"0" & TYPE_4 & I_SEND when X"655",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"656",
            X"020" when X"657",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"658",
            X"004" when X"659",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"65A",
            X"020" when X"65B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"65C",
            X"005" when X"65D",
            X"0" & TYPE_4 & I_SEND when X"65E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"65F",
            X"04F" when X"660",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"661",
            X"004" when X"662",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"663",
            X"04B" when X"664",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"665",
            X"005" when X"666",
            X"0" & TYPE_4 & I_SEND when X"667",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"668",
            X"044" when X"669",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"66A",
            X"009" when X"66B",
            X"0" & TYPE_2 & JMP_UNCOND when X"66C",
            X"880" when X"66D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"66E",
            X"001" when X"66F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"670",
            X"038" when X"671",
            X"0" & TYPE_1 & ALU_CMPE when X"672",
            X"0" & TYPE_2 & JMP_COND when X"673",
            X"677" when X"674",
            X"0" & TYPE_2 & JMP_UNCOND when X"675",
            X"6E0" when X"676",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"677",
            X"044" when X"678",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"679",
            X"005" when X"67A",
            X"0" & TYPE_1 & ALU_CMPL when X"67B",
            X"0" & TYPE_2 & JMP_COND when X"67C",
            X"680" when X"67D",
            X"0" & TYPE_2 & JMP_UNCOND when X"67E",
            X"68B" when X"67F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"680",
            X"045" when X"681",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"682",
            X"004" when X"683",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"684",
            X"052" when X"685",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"686",
            X"005" when X"687",
            X"0" & TYPE_4 & I_SEND when X"688",
            X"0" & TYPE_2 & JMP_UNCOND when X"689",
            X"880" when X"68A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"68B",
            X"044" when X"68C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"68D",
            X"008" when X"68E",
            X"0" & TYPE_1 & ALU_CMPG when X"68F",
            X"0" & TYPE_2 & JMP_COND when X"690",
            X"694" when X"691",
            X"0" & TYPE_2 & JMP_UNCOND when X"692",
            X"69F" when X"693",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"694",
            X"045" when X"695",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"696",
            X"004" when X"697",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"698",
            X"052" when X"699",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"69A",
            X"005" when X"69B",
            X"0" & TYPE_4 & I_SEND when X"69C",
            X"0" & TYPE_2 & JMP_UNCOND when X"69D",
            X"880" when X"69E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"69F",
            X"04E" when X"6A0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6A1",
            X"004" when X"6A2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6A3",
            X"05F" when X"6A4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6A5",
            X"005" when X"6A6",
            X"0" & TYPE_4 & I_SEND when X"6A7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6A8",
            X"042" when X"6A9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6AA",
            X"004" when X"6AB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6AC",
            X"049" when X"6AD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6AE",
            X"005" when X"6AF",
            X"0" & TYPE_4 & I_SEND when X"6B0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6B1",
            X"054" when X"6B2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6B3",
            X"004" when X"6B4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6B5",
            X"053" when X"6B6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6B7",
            X"005" when X"6B8",
            X"0" & TYPE_4 & I_SEND when X"6B9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6BA",
            X"03A" when X"6BB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6BC",
            X"004" when X"6BD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6BE",
            X"020" when X"6BF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6C0",
            X"005" when X"6C1",
            X"0" & TYPE_4 & I_SEND when X"6C2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"6C3",
            X"002" when X"6C4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"6C5",
            X"030" when X"6C6",
            X"0" & TYPE_1 & ALU_SUB when X"6C7",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"6C8",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"6C9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6CA",
            X"004" when X"6CB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6CC",
            X"020" when X"6CD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6CE",
            X"005" when X"6CF",
            X"0" & TYPE_4 & I_SEND when X"6D0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6D1",
            X"04F" when X"6D2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6D3",
            X"004" when X"6D4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6D5",
            X"04B" when X"6D6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6D7",
            X"005" when X"6D8",
            X"0" & TYPE_4 & I_SEND when X"6D9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"6DA",
            X"044" when X"6DB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6DC",
            X"008" when X"6DD",
            X"0" & TYPE_2 & JMP_UNCOND when X"6DE",
            X"880" when X"6DF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"6E0",
            X"001" when X"6E1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"6E2",
            X"037" when X"6E3",
            X"0" & TYPE_1 & ALU_CMPE when X"6E4",
            X"0" & TYPE_2 & JMP_COND when X"6E5",
            X"6E9" when X"6E6",
            X"0" & TYPE_2 & JMP_UNCOND when X"6E7",
            X"77A" when X"6E8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"6E9",
            X"044" when X"6EA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"6EB",
            X"002" when X"6EC",
            X"0" & TYPE_1 & ALU_CMPL when X"6ED",
            X"0" & TYPE_2 & JMP_COND when X"6EE",
            X"6F2" when X"6EF",
            X"0" & TYPE_2 & JMP_UNCOND when X"6F0",
            X"6FD" when X"6F1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6F2",
            X"045" when X"6F3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6F4",
            X"004" when X"6F5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"6F6",
            X"052" when X"6F7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"6F8",
            X"005" when X"6F9",
            X"0" & TYPE_4 & I_SEND when X"6FA",
            X"0" & TYPE_2 & JMP_UNCOND when X"6FB",
            X"880" when X"6FC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"6FD",
            X"044" when X"6FE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"6FF",
            X"004" when X"700",
            X"0" & TYPE_1 & ALU_CMPG when X"701",
            X"0" & TYPE_2 & JMP_COND when X"702",
            X"706" when X"703",
            X"0" & TYPE_2 & JMP_UNCOND when X"704",
            X"711" when X"705",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"706",
            X"045" when X"707",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"708",
            X"004" when X"709",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"70A",
            X"052" when X"70B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"70C",
            X"005" when X"70D",
            X"0" & TYPE_4 & I_SEND when X"70E",
            X"0" & TYPE_2 & JMP_UNCOND when X"70F",
            X"880" when X"710",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"711",
            X"053" when X"712",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"713",
            X"004" when X"714",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"715",
            X"054" when X"716",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"717",
            X"005" when X"718",
            X"0" & TYPE_4 & I_SEND when X"719",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"71A",
            X"04F" when X"71B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"71C",
            X"004" when X"71D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"71E",
            X"050" when X"71F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"720",
            X"005" when X"721",
            X"0" & TYPE_4 & I_SEND when X"722",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"723",
            X"03A" when X"724",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"725",
            X"004" when X"726",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"727",
            X"020" when X"728",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"729",
            X"005" when X"72A",
            X"0" & TYPE_4 & I_SEND when X"72B",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"72C",
            X"002" when X"72D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"72E",
            X"032" when X"72F",
            X"0" & TYPE_1 & ALU_CMPE when X"730",
            X"0" & TYPE_2 & JMP_COND when X"731",
            X"735" when X"732",
            X"0" & TYPE_2 & JMP_UNCOND when X"733",
            X"73E" when X"734",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"735",
            X"031" when X"736",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"737",
            X"004" when X"738",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"739",
            X"020" when X"73A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"73B",
            X"005" when X"73C",
            X"0" & TYPE_4 & I_SEND when X"73D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"73E",
            X"002" when X"73F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"740",
            X"033" when X"741",
            X"0" & TYPE_1 & ALU_CMPE when X"742",
            X"0" & TYPE_2 & JMP_COND when X"743",
            X"747" when X"744",
            X"0" & TYPE_2 & JMP_UNCOND when X"745",
            X"759" when X"746",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"747",
            X"031" when X"748",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"749",
            X"004" when X"74A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"74B",
            X"02E" when X"74C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"74D",
            X"005" when X"74E",
            X"0" & TYPE_4 & I_SEND when X"74F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"750",
            X"035" when X"751",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"752",
            X"004" when X"753",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"754",
            X"020" when X"755",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"756",
            X"005" when X"757",
            X"0" & TYPE_4 & I_SEND when X"758",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"759",
            X"002" when X"75A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"75B",
            X"034" when X"75C",
            X"0" & TYPE_1 & ALU_CMPE when X"75D",
            X"0" & TYPE_2 & JMP_COND when X"75E",
            X"762" when X"75F",
            X"0" & TYPE_2 & JMP_UNCOND when X"760",
            X"76B" when X"761",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"762",
            X"032" when X"763",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"764",
            X"004" when X"765",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"766",
            X"020" when X"767",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"768",
            X"005" when X"769",
            X"0" & TYPE_4 & I_SEND when X"76A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"76B",
            X"04F" when X"76C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"76D",
            X"004" when X"76E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"76F",
            X"04B" when X"770",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"771",
            X"005" when X"772",
            X"0" & TYPE_4 & I_SEND when X"773",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"774",
            X"044" when X"775",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"776",
            X"007" when X"777",
            X"0" & TYPE_2 & JMP_UNCOND when X"778",
            X"880" when X"779",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"77A",
            X"001" when X"77B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"77C",
            X"036" when X"77D",
            X"0" & TYPE_1 & ALU_CMPE when X"77E",
            X"0" & TYPE_2 & JMP_COND when X"77F",
            X"783" when X"780",
            X"0" & TYPE_2 & JMP_UNCOND when X"781",
            X"875" when X"782",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"783",
            X"044" when X"784",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"785",
            X"004" when X"786",
            X"0" & TYPE_1 & ALU_CMPG when X"787",
            X"0" & TYPE_2 & JMP_COND when X"788",
            X"78C" when X"789",
            X"0" & TYPE_2 & JMP_UNCOND when X"78A",
            X"797" when X"78B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"78C",
            X"045" when X"78D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"78E",
            X"004" when X"78F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"790",
            X"052" when X"791",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"792",
            X"005" when X"793",
            X"0" & TYPE_4 & I_SEND when X"794",
            X"0" & TYPE_2 & JMP_UNCOND when X"795",
            X"880" when X"796",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"797",
            X"050" when X"798",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"799",
            X"004" when X"79A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"79B",
            X"041" when X"79C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"79D",
            X"005" when X"79E",
            X"0" & TYPE_4 & I_SEND when X"79F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7A0",
            X"052" when X"7A1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7A2",
            X"004" when X"7A3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7A4",
            X"049" when X"7A5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7A6",
            X"005" when X"7A7",
            X"0" & TYPE_4 & I_SEND when X"7A8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7A9",
            X"054" when X"7AA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7AB",
            X"004" when X"7AC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7AD",
            X"059" when X"7AE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7AF",
            X"005" when X"7B0",
            X"0" & TYPE_4 & I_SEND when X"7B1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7B2",
            X"03A" when X"7B3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7B4",
            X"004" when X"7B5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7B6",
            X"020" when X"7B7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7B8",
            X"005" when X"7B9",
            X"0" & TYPE_4 & I_SEND when X"7BA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"7BB",
            X"002" when X"7BC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"7BD",
            X"030" when X"7BE",
            X"0" & TYPE_1 & ALU_CMPE when X"7BF",
            X"0" & TYPE_2 & JMP_COND when X"7C0",
            X"7C4" when X"7C1",
            X"0" & TYPE_2 & JMP_UNCOND when X"7C2",
            X"7DF" when X"7C3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7C4",
            X"045" when X"7C5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7C6",
            X"004" when X"7C7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7C8",
            X"056" when X"7C9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7CA",
            X"005" when X"7CB",
            X"0" & TYPE_4 & I_SEND when X"7CC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7CD",
            X"045" when X"7CE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7CF",
            X"004" when X"7D0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7D1",
            X"04E" when X"7D2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7D3",
            X"005" when X"7D4",
            X"0" & TYPE_4 & I_SEND when X"7D5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7D6",
            X"020" when X"7D7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7D8",
            X"004" when X"7D9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7DA",
            X"020" when X"7DB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7DC",
            X"005" when X"7DD",
            X"0" & TYPE_4 & I_SEND when X"7DE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"7DF",
            X"002" when X"7E0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"7E1",
            X"031" when X"7E2",
            X"0" & TYPE_1 & ALU_CMPE when X"7E3",
            X"0" & TYPE_2 & JMP_COND when X"7E4",
            X"7E8" when X"7E5",
            X"0" & TYPE_2 & JMP_UNCOND when X"7E6",
            X"7FA" when X"7E7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7E8",
            X"04F" when X"7E9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7EA",
            X"004" when X"7EB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7EC",
            X"044" when X"7ED",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7EE",
            X"005" when X"7EF",
            X"0" & TYPE_4 & I_SEND when X"7F0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7F1",
            X"044" when X"7F2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7F3",
            X"004" when X"7F4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"7F5",
            X"020" when X"7F6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"7F7",
            X"005" when X"7F8",
            X"0" & TYPE_4 & I_SEND when X"7F9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"7FA",
            X"002" when X"7FB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"7FC",
            X"032" when X"7FD",
            X"0" & TYPE_1 & ALU_CMPE when X"7FE",
            X"0" & TYPE_2 & JMP_COND when X"7FF",
            X"803" when X"800",
            X"0" & TYPE_2 & JMP_UNCOND when X"801",
            X"81E" when X"802",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"803",
            X"04D" when X"804",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"805",
            X"004" when X"806",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"807",
            X"041" when X"808",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"809",
            X"005" when X"80A",
            X"0" & TYPE_4 & I_SEND when X"80B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"80C",
            X"052" when X"80D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"80E",
            X"004" when X"80F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"810",
            X"04B" when X"811",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"812",
            X"005" when X"813",
            X"0" & TYPE_4 & I_SEND when X"814",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"815",
            X"020" when X"816",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"817",
            X"004" when X"818",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"819",
            X"020" when X"81A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"81B",
            X"005" when X"81C",
            X"0" & TYPE_4 & I_SEND when X"81D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"81E",
            X"002" when X"81F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"820",
            X"033" when X"821",
            X"0" & TYPE_1 & ALU_CMPE when X"822",
            X"0" & TYPE_2 & JMP_COND when X"823",
            X"827" when X"824",
            X"0" & TYPE_2 & JMP_UNCOND when X"825",
            X"842" when X"826",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"827",
            X"053" when X"828",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"829",
            X"004" when X"82A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"82B",
            X"050" when X"82C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"82D",
            X"005" when X"82E",
            X"0" & TYPE_4 & I_SEND when X"82F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"830",
            X"041" when X"831",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"832",
            X"004" when X"833",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"834",
            X"043" when X"835",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"836",
            X"005" when X"837",
            X"0" & TYPE_4 & I_SEND when X"838",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"839",
            X"045" when X"83A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"83B",
            X"004" when X"83C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"83D",
            X"020" when X"83E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"83F",
            X"005" when X"840",
            X"0" & TYPE_4 & I_SEND when X"841",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"842",
            X"002" when X"843",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"844",
            X"034" when X"845",
            X"0" & TYPE_1 & ALU_CMPE when X"846",
            X"0" & TYPE_2 & JMP_COND when X"847",
            X"84B" when X"848",
            X"0" & TYPE_2 & JMP_UNCOND when X"849",
            X"866" when X"84A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"84B",
            X"04E" when X"84C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"84D",
            X"004" when X"84E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"84F",
            X"04F" when X"850",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"851",
            X"005" when X"852",
            X"0" & TYPE_4 & I_SEND when X"853",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"854",
            X"04E" when X"855",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"856",
            X"004" when X"857",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"858",
            X"045" when X"859",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"85A",
            X"005" when X"85B",
            X"0" & TYPE_4 & I_SEND when X"85C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"85D",
            X"020" when X"85E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"85F",
            X"004" when X"860",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"861",
            X"020" when X"862",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"863",
            X"005" when X"864",
            X"0" & TYPE_4 & I_SEND when X"865",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"866",
            X"04F" when X"867",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"868",
            X"004" when X"869",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"86A",
            X"04B" when X"86B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"86C",
            X"005" when X"86D",
            X"0" & TYPE_4 & I_SEND when X"86E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"86F",
            X"044" when X"870",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"871",
            X"050" when X"872",
            X"0" & TYPE_2 & JMP_UNCOND when X"873",
            X"880" when X"874",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"875",
            X"045" when X"876",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"877",
            X"004" when X"878",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"879",
            X"052" when X"87A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"87B",
            X"005" when X"87C",
            X"0" & TYPE_4 & I_SEND when X"87D",
            X"0" & TYPE_2 & JMP_UNCOND when X"87E",
            X"880" when X"87F",
            X"0" & TYPE_4 & I_RETI when X"880",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"881",
            X"000" when X"882",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"883",
            X"04F" when X"884",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"885",
            X"004" when X"886",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"887",
            X"050" when X"888",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"889",
            X"002" when X"88A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"88B",
            X"007" when X"88C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"88D",
            X"008" when X"88E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"88F",
            X"008" when X"890",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"891",
            X"008" when X"892",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"893",
            X"009" when X"894",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"895",
            X"010" when X"896",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"897",
            X"031" when X"898",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"899",
            X"000" when X"89A",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"89B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"89C",
            X"000" when X"89D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"89E",
            X"020" when X"89F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8A0",
            X"000" when X"8A1",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"8A2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8A3",
            X"000" when X"8A4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"8A5",
            X"010" when X"8A6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8A7",
            X"000" when X"8A8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8A9",
            X"003" when X"8AA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8AB",
            X"04C" when X"8AC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8AD",
            X"051" when X"8AE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8AF",
            X"000" when X"8B0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8B1",
            X"052" when X"8B2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8B3",
            X"051" when X"8B4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8B5",
            X"053" when X"8B6",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8B7",
            X"051" when X"8B8",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8B9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8BA",
            X"008" when X"8BB",
            X"0" & TYPE_1 & ALU_CMPL when X"8BC",
            X"0" & TYPE_2 & JMP_COND when X"8BD",
            X"8E1" when X"8BE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8BF",
            X"051" when X"8C0",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8C1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8C2",
            X"010" when X"8C3",
            X"0" & TYPE_1 & ALU_CMPL when X"8C4",
            X"0" & TYPE_2 & JMP_COND when X"8C5",
            X"8D5" when X"8C6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8C7",
            X"002" when X"8C8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8C9",
            X"052" when X"8CA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8CB",
            X"051" when X"8CC",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8CD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8CE",
            X"010" when X"8CF",
            X"0" & TYPE_1 & ALU_SUB when X"8D0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8D1",
            X"053" when X"8D2",
            X"0" & TYPE_2 & JMP_UNCOND when X"8D3",
            X"8E1" when X"8D4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8D5",
            X"001" when X"8D6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8D7",
            X"052" when X"8D8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8D9",
            X"051" when X"8DA",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8DB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8DC",
            X"008" when X"8DD",
            X"0" & TYPE_1 & ALU_SUB when X"8DE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8DF",
            X"053" when X"8E0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"8E1",
            X"001" when X"8E2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8E3",
            X"054" when X"8E4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8E5",
            X"053" when X"8E6",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8E7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8E8",
            X"000" when X"8E9",
            X"0" & TYPE_1 & ALU_CMPE when X"8EA",
            X"0" & TYPE_2 & JMP_COND when X"8EB",
            X"900" when X"8EC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8ED",
            X"054" when X"8EE",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8EF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8F0",
            X"000" when X"8F1",
            X"0" & TYPE_1 & ALU_ADD when X"8F2",
            X"0" & TYPE_1 & ALU_SHIFTL when X"8F3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8F4",
            X"054" when X"8F5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"8F6",
            X"053" when X"8F7",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"8F8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"8F9",
            X"001" when X"8FA",
            X"0" & TYPE_1 & ALU_SUB when X"8FB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"8FC",
            X"053" when X"8FD",
            X"0" & TYPE_2 & JMP_UNCOND when X"8FE",
            X"8E5" when X"8FF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"900",
            X"052" when X"901",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"902",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"903",
            X"01B" when X"904",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"905",
            X"041" when X"906",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"907",
            X"054" when X"908",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_B when X"909",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"90A",
            X"041" when X"90B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"90C",
            X"0" & TYPE_1 & ALU_OR when X"90D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"90E",
            X"041" when X"90F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"910",
            X"052" when X"911",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"912",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"913",
            X"041" when X"914",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"915",
            X"01B" when X"916",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"917",
            X"053" when X"918",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"919",
            X"004" when X"91A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"91B",
            X"059" when X"91C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"91D",
            X"005" when X"91E",
            X"0" & TYPE_4 & I_SEND when X"91F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"920",
            X"053" when X"921",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"922",
            X"004" when X"923",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"924",
            X"054" when X"925",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"926",
            X"005" when X"927",
            X"0" & TYPE_4 & I_SEND when X"928",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"929",
            X"045" when X"92A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"92B",
            X"004" when X"92C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"92D",
            X"04D" when X"92E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"92F",
            X"005" when X"930",
            X"0" & TYPE_4 & I_SEND when X"931",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"932",
            X"020" when X"933",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"934",
            X"004" when X"935",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"936",
            X"052" when X"937",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"938",
            X"005" when X"939",
            X"0" & TYPE_4 & I_SEND when X"93A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"93B",
            X"045" when X"93C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"93D",
            X"004" when X"93E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"93F",
            X"041" when X"940",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"941",
            X"005" when X"942",
            X"0" & TYPE_4 & I_SEND when X"943",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"944",
            X"044" when X"945",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"946",
            X"004" when X"947",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"948",
            X"059" when X"949",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"94A",
            X"005" when X"94B",
            X"0" & TYPE_4 & I_SEND when X"94C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"94D",
            X"00A" when X"94E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"94F",
            X"004" when X"950",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"951",
            X"020" when X"952",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"953",
            X"005" when X"954",
            X"0" & TYPE_4 & I_SEND when X"955",
            X"0" & TYPE_2 & JMP_UNCOND when X"956",
            X"958" when X"957",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"958",
            X"019" when X"959",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"95A",
            X"000" when X"95B",
            X"0" & TYPE_1 & ALU_ADD when X"95C",
            X"0" & TYPE_1 & ALU_SHIFTR when X"95D",
            X"0" & TYPE_1 & ALU_SHIFTR when X"95E",
            X"0" & TYPE_1 & ALU_SHIFTR when X"95F",
            X"0" & TYPE_1 & ALU_SHIFTR when X"960",
            X"0" & TYPE_1 & ALU_SHIFTR when X"961",
            X"0" & TYPE_1 & ALU_SHIFTR when X"962",
            X"0" & TYPE_1 & ALU_SHIFTR when X"963",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"964",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"965",
            X"001" when X"966",
            X"0" & TYPE_1 & ALU_AND when X"967",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"968",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"969",
            X"001" when X"96A",
            X"0" & TYPE_1 & ALU_CMPE when X"96B",
            X"0" & TYPE_2 & JMP_COND when X"96C",
            X"970" when X"96D",
            X"0" & TYPE_2 & JMP_UNCOND when X"96E",
            X"9F5" when X"96F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"970",
            X"047" when X"971",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"972",
            X"000" when X"973",
            X"0" & TYPE_1 & ALU_CMPE when X"974",
            X"0" & TYPE_2 & JMP_COND when X"975",
            X"979" when X"976",
            X"0" & TYPE_2 & JMP_UNCOND when X"977",
            X"9F5" when X"978",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"979",
            X"001" when X"97A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"97B",
            X"047" when X"97C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"97D",
            X"042" when X"97E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"97F",
            X"004" when X"980",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"981",
            X"06F" when X"982",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"983",
            X"005" when X"984",
            X"0" & TYPE_4 & I_SEND when X"985",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"986",
            X"074" when X"987",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"988",
            X"004" when X"989",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"98A",
            X"06F" when X"98B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"98C",
            X"005" when X"98D",
            X"0" & TYPE_4 & I_SEND when X"98E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"98F",
            X"06E" when X"990",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"991",
            X"004" when X"992",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"993",
            X"020" when X"994",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"995",
            X"005" when X"996",
            X"0" & TYPE_4 & I_SEND when X"997",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"998",
            X"055" when X"999",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"99A",
            X"004" when X"99B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"99C",
            X"050" when X"99D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"99E",
            X"005" when X"99F",
            X"0" & TYPE_4 & I_SEND when X"9A0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9A1",
            X"020" when X"9A2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9A3",
            X"004" when X"9A4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9A5",
            X"070" when X"9A6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9A7",
            X"005" when X"9A8",
            X"0" & TYPE_4 & I_SEND when X"9A9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9AA",
            X"075" when X"9AB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9AC",
            X"004" when X"9AD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9AE",
            X"06C" when X"9AF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9B0",
            X"005" when X"9B1",
            X"0" & TYPE_4 & I_SEND when X"9B2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9B3",
            X"073" when X"9B4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9B5",
            X"004" when X"9B6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9B7",
            X"061" when X"9B8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9B9",
            X"005" when X"9BA",
            X"0" & TYPE_4 & I_SEND when X"9BB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9BC",
            X"064" when X"9BD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9BE",
            X"004" when X"9BF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9C0",
            X"06F" when X"9C1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9C2",
            X"005" when X"9C3",
            X"0" & TYPE_4 & I_SEND when X"9C4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9C5",
            X"00A" when X"9C6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9C7",
            X"004" when X"9C8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"9C9",
            X"020" when X"9CA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9CB",
            X"005" when X"9CC",
            X"0" & TYPE_4 & I_SEND when X"9CD",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9CE",
            X"031" when X"9CF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9D0",
            X"029" when X"9D1",
            X"0" & TYPE_1 & ALU_CMPL when X"9D2",
            X"0" & TYPE_2 & JMP_COND when X"9D3",
            X"9D7" when X"9D4",
            X"0" & TYPE_2 & JMP_UNCOND when X"9D5",
            X"9F5" when X"9D6",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9D7",
            X"031" when X"9D8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9D9",
            X"001" when X"9DA",
            X"0" & TYPE_1 & ALU_ADD when X"9DB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9DC",
            X"031" when X"9DD",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9DE",
            X"031" when X"9DF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9E0",
            X"00F" when X"9E1",
            X"0" & TYPE_1 & ALU_AND when X"9E2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9E3",
            X"046" when X"9E4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9E5",
            X"046" when X"9E6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9E7",
            X"009" when X"9E8",
            X"0" & TYPE_1 & ALU_CMPG when X"9E9",
            X"0" & TYPE_2 & JMP_COND when X"9EA",
            X"9EE" when X"9EB",
            X"0" & TYPE_2 & JMP_UNCOND when X"9EC",
            X"9F5" when X"9ED",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9EE",
            X"031" when X"9EF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9F0",
            X"006" when X"9F1",
            X"0" & TYPE_1 & ALU_ADD when X"9F2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"9F3",
            X"031" when X"9F4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"9F5",
            X"019" when X"9F6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"9F7",
            X"000" when X"9F8",
            X"0" & TYPE_1 & ALU_ADD when X"9F9",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FA",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FB",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FC",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FD",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FE",
            X"0" & TYPE_1 & ALU_SHIFTR when X"9FF",
            X"0" & TYPE_1 & ALU_SHIFTR when X"A00",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"A01",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A02",
            X"001" when X"A03",
            X"0" & TYPE_1 & ALU_AND when X"A04",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"A05",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A06",
            X"000" when X"A07",
            X"0" & TYPE_1 & ALU_CMPE when X"A08",
            X"0" & TYPE_2 & JMP_COND when X"A09",
            X"A0D" when X"A0A",
            X"0" & TYPE_2 & JMP_UNCOND when X"A0B",
            X"A11" when X"A0C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A0D",
            X"000" when X"A0E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A0F",
            X"047" when X"A10",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"A11",
            X"01A" when X"A12",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A13",
            X"000" when X"A14",
            X"0" & TYPE_1 & ALU_ADD when X"A15",
            X"0" & TYPE_1 & ALU_SHIFTR when X"A16",
            X"0" & TYPE_1 & ALU_SHIFTR when X"A17",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"A18",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A19",
            X"001" when X"A1A",
            X"0" & TYPE_1 & ALU_AND when X"A1B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"A1C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A1D",
            X"001" when X"A1E",
            X"0" & TYPE_1 & ALU_CMPE when X"A1F",
            X"0" & TYPE_2 & JMP_COND when X"A20",
            X"A24" when X"A21",
            X"0" & TYPE_2 & JMP_UNCOND when X"A22",
            X"AB2" when X"A23",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"A24",
            X"048" when X"A25",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A26",
            X"000" when X"A27",
            X"0" & TYPE_1 & ALU_CMPE when X"A28",
            X"0" & TYPE_2 & JMP_COND when X"A29",
            X"A2D" when X"A2A",
            X"0" & TYPE_2 & JMP_UNCOND when X"A2B",
            X"AB2" when X"A2C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A2D",
            X"001" when X"A2E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A2F",
            X"048" when X"A30",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A31",
            X"042" when X"A32",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A33",
            X"004" when X"A34",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A35",
            X"06F" when X"A36",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A37",
            X"005" when X"A38",
            X"0" & TYPE_4 & I_SEND when X"A39",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A3A",
            X"074" when X"A3B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A3C",
            X"004" when X"A3D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A3E",
            X"06F" when X"A3F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A40",
            X"005" when X"A41",
            X"0" & TYPE_4 & I_SEND when X"A42",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A43",
            X"06E" when X"A44",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A45",
            X"004" when X"A46",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A47",
            X"020" when X"A48",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A49",
            X"005" when X"A4A",
            X"0" & TYPE_4 & I_SEND when X"A4B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A4C",
            X"044" when X"A4D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A4E",
            X"004" when X"A4F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A50",
            X"04F" when X"A51",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A52",
            X"005" when X"A53",
            X"0" & TYPE_4 & I_SEND when X"A54",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A55",
            X"057" when X"A56",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A57",
            X"004" when X"A58",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A59",
            X"04E" when X"A5A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A5B",
            X"005" when X"A5C",
            X"0" & TYPE_4 & I_SEND when X"A5D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A5E",
            X"020" when X"A5F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A60",
            X"004" when X"A61",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A62",
            X"070" when X"A63",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A64",
            X"005" when X"A65",
            X"0" & TYPE_4 & I_SEND when X"A66",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A67",
            X"075" when X"A68",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A69",
            X"004" when X"A6A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A6B",
            X"06C" when X"A6C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A6D",
            X"005" when X"A6E",
            X"0" & TYPE_4 & I_SEND when X"A6F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A70",
            X"073" when X"A71",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A72",
            X"004" when X"A73",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A74",
            X"061" when X"A75",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A76",
            X"005" when X"A77",
            X"0" & TYPE_4 & I_SEND when X"A78",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A79",
            X"064" when X"A7A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A7B",
            X"004" when X"A7C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A7D",
            X"06F" when X"A7E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A7F",
            X"005" when X"A80",
            X"0" & TYPE_4 & I_SEND when X"A81",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A82",
            X"00A" when X"A83",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A84",
            X"004" when X"A85",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"A86",
            X"020" when X"A87",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A88",
            X"005" when X"A89",
            X"0" & TYPE_4 & I_SEND when X"A8A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"A8B",
            X"031" when X"A8C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A8D",
            X"000" when X"A8E",
            X"0" & TYPE_1 & ALU_CMPG when X"A8F",
            X"0" & TYPE_2 & JMP_COND when X"A90",
            X"A94" when X"A91",
            X"0" & TYPE_2 & JMP_UNCOND when X"A92",
            X"AB2" when X"A93",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"A94",
            X"031" when X"A95",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A96",
            X"001" when X"A97",
            X"0" & TYPE_1 & ALU_SUB when X"A98",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"A99",
            X"031" when X"A9A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"A9B",
            X"031" when X"A9C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"A9D",
            X"00F" when X"A9E",
            X"0" & TYPE_1 & ALU_AND when X"A9F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AA0",
            X"046" when X"AA1",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"AA2",
            X"046" when X"AA3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"AA4",
            X"009" when X"AA5",
            X"0" & TYPE_1 & ALU_CMPG when X"AA6",
            X"0" & TYPE_2 & JMP_COND when X"AA7",
            X"AAB" when X"AA8",
            X"0" & TYPE_2 & JMP_UNCOND when X"AA9",
            X"AB2" when X"AAA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"AAB",
            X"031" when X"AAC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"AAD",
            X"006" when X"AAE",
            X"0" & TYPE_1 & ALU_SUB when X"AAF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AB0",
            X"031" when X"AB1",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"AB2",
            X"01A" when X"AB3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"AB4",
            X"000" when X"AB5",
            X"0" & TYPE_1 & ALU_ADD when X"AB6",
            X"0" & TYPE_1 & ALU_SHIFTR when X"AB7",
            X"0" & TYPE_1 & ALU_SHIFTR when X"AB8",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"AB9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ABA",
            X"001" when X"ABB",
            X"0" & TYPE_1 & ALU_AND when X"ABC",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"ABD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ABE",
            X"000" when X"ABF",
            X"0" & TYPE_1 & ALU_CMPE when X"AC0",
            X"0" & TYPE_2 & JMP_COND when X"AC1",
            X"AC5" when X"AC2",
            X"0" & TYPE_2 & JMP_UNCOND when X"AC3",
            X"AC9" when X"AC4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AC5",
            X"000" when X"AC6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AC7",
            X"048" when X"AC8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"AC9",
            X"01A" when X"ACA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ACB",
            X"000" when X"ACC",
            X"0" & TYPE_1 & ALU_ADD when X"ACD",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"ACE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ACF",
            X"001" when X"AD0",
            X"0" & TYPE_1 & ALU_AND when X"AD1",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"AD2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"AD3",
            X"001" when X"AD4",
            X"0" & TYPE_1 & ALU_CMPE when X"AD5",
            X"0" & TYPE_2 & JMP_COND when X"AD6",
            X"ADA" when X"AD7",
            X"0" & TYPE_2 & JMP_UNCOND when X"AD8",
            X"C2D" when X"AD9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"ADA",
            X"049" when X"ADB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ADC",
            X"000" when X"ADD",
            X"0" & TYPE_1 & ALU_CMPE when X"ADE",
            X"0" & TYPE_2 & JMP_COND when X"ADF",
            X"AE3" when X"AE0",
            X"0" & TYPE_2 & JMP_UNCOND when X"AE1",
            X"C2D" when X"AE2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AE3",
            X"001" when X"AE4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AE5",
            X"049" when X"AE6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AE7",
            X"042" when X"AE8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AE9",
            X"004" when X"AEA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AEB",
            X"06F" when X"AEC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AED",
            X"005" when X"AEE",
            X"0" & TYPE_4 & I_SEND when X"AEF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AF0",
            X"074" when X"AF1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AF2",
            X"004" when X"AF3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AF4",
            X"06F" when X"AF5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AF6",
            X"005" when X"AF7",
            X"0" & TYPE_4 & I_SEND when X"AF8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AF9",
            X"06E" when X"AFA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AFB",
            X"004" when X"AFC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"AFD",
            X"020" when X"AFE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"AFF",
            X"005" when X"B00",
            X"0" & TYPE_4 & I_SEND when X"B01",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B02",
            X"04C" when X"B03",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B04",
            X"004" when X"B05",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B06",
            X"045" when X"B07",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B08",
            X"005" when X"B09",
            X"0" & TYPE_4 & I_SEND when X"B0A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B0B",
            X"046" when X"B0C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B0D",
            X"004" when X"B0E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B0F",
            X"054" when X"B10",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B11",
            X"005" when X"B12",
            X"0" & TYPE_4 & I_SEND when X"B13",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B14",
            X"020" when X"B15",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B16",
            X"004" when X"B17",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B18",
            X"070" when X"B19",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B1A",
            X"005" when X"B1B",
            X"0" & TYPE_4 & I_SEND when X"B1C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B1D",
            X"075" when X"B1E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B1F",
            X"004" when X"B20",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B21",
            X"06C" when X"B22",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B23",
            X"005" when X"B24",
            X"0" & TYPE_4 & I_SEND when X"B25",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B26",
            X"073" when X"B27",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B28",
            X"004" when X"B29",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B2A",
            X"061" when X"B2B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B2C",
            X"005" when X"B2D",
            X"0" & TYPE_4 & I_SEND when X"B2E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B2F",
            X"064" when X"B30",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B31",
            X"004" when X"B32",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B33",
            X"06F" when X"B34",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B35",
            X"005" when X"B36",
            X"0" & TYPE_4 & I_SEND when X"B37",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B38",
            X"00A" when X"B39",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B3A",
            X"004" when X"B3B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B3C",
            X"020" when X"B3D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B3E",
            X"005" when X"B3F",
            X"0" & TYPE_4 & I_SEND when X"B40",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"B41",
            X"04C" when X"B42",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B43",
            X"007" when X"B44",
            X"0" & TYPE_1 & ALU_CMPL when X"B45",
            X"0" & TYPE_2 & JMP_COND when X"B46",
            X"B4A" when X"B47",
            X"0" & TYPE_2 & JMP_UNCOND when X"B48",
            X"C2D" when X"B49",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B4A",
            X"04C" when X"B4B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B4C",
            X"051" when X"B4D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B4E",
            X"000" when X"B4F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B50",
            X"052" when X"B51",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B52",
            X"051" when X"B53",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B54",
            X"053" when X"B55",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B56",
            X"051" when X"B57",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B58",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B59",
            X"008" when X"B5A",
            X"0" & TYPE_1 & ALU_CMPL when X"B5B",
            X"0" & TYPE_2 & JMP_COND when X"B5C",
            X"B80" when X"B5D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B5E",
            X"051" when X"B5F",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B60",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B61",
            X"010" when X"B62",
            X"0" & TYPE_1 & ALU_CMPL when X"B63",
            X"0" & TYPE_2 & JMP_COND when X"B64",
            X"B74" when X"B65",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B66",
            X"002" when X"B67",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B68",
            X"052" when X"B69",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B6A",
            X"051" when X"B6B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B6C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B6D",
            X"010" when X"B6E",
            X"0" & TYPE_1 & ALU_SUB when X"B6F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B70",
            X"053" when X"B71",
            X"0" & TYPE_2 & JMP_UNCOND when X"B72",
            X"B80" when X"B73",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B74",
            X"001" when X"B75",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B76",
            X"052" when X"B77",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B78",
            X"051" when X"B79",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B7A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B7B",
            X"008" when X"B7C",
            X"0" & TYPE_1 & ALU_SUB when X"B7D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B7E",
            X"053" when X"B7F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"B80",
            X"001" when X"B81",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B82",
            X"054" when X"B83",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B84",
            X"053" when X"B85",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B86",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B87",
            X"000" when X"B88",
            X"0" & TYPE_1 & ALU_CMPE when X"B89",
            X"0" & TYPE_2 & JMP_COND when X"B8A",
            X"B9F" when X"B8B",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B8C",
            X"054" when X"B8D",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B8E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B8F",
            X"000" when X"B90",
            X"0" & TYPE_1 & ALU_ADD when X"B91",
            X"0" & TYPE_1 & ALU_SHIFTL when X"B92",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B93",
            X"054" when X"B94",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B95",
            X"053" when X"B96",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"B97",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"B98",
            X"001" when X"B99",
            X"0" & TYPE_1 & ALU_SUB when X"B9A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"B9B",
            X"053" when X"B9C",
            X"0" & TYPE_2 & JMP_UNCOND when X"B9D",
            X"B84" when X"B9E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"B9F",
            X"052" when X"BA0",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"BA1",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"BA2",
            X"01B" when X"BA3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BA4",
            X"041" when X"BA5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BA6",
            X"054" when X"BA7",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BA8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BA9",
            X"0FF" when X"BAA",
            X"0" & TYPE_1 & ALU_XOR when X"BAB",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_B when X"BAC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BAD",
            X"041" when X"BAE",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BAF",
            X"0" & TYPE_1 & ALU_AND when X"BB0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BB1",
            X"041" when X"BB2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BB3",
            X"052" when X"BB4",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"BB5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BB6",
            X"041" when X"BB7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"BB8",
            X"01B" when X"BB9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"BBA",
            X"04C" when X"BBB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BBC",
            X"001" when X"BBD",
            X"0" & TYPE_1 & ALU_ADD when X"BBE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BBF",
            X"04C" when X"BC0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BC1",
            X"04C" when X"BC2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BC3",
            X"051" when X"BC4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"BC5",
            X"000" when X"BC6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BC7",
            X"052" when X"BC8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BC9",
            X"051" when X"BCA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BCB",
            X"053" when X"BCC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BCD",
            X"051" when X"BCE",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BCF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BD0",
            X"008" when X"BD1",
            X"0" & TYPE_1 & ALU_CMPL when X"BD2",
            X"0" & TYPE_2 & JMP_COND when X"BD3",
            X"BF7" when X"BD4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BD5",
            X"051" when X"BD6",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BD7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BD8",
            X"010" when X"BD9",
            X"0" & TYPE_1 & ALU_CMPL when X"BDA",
            X"0" & TYPE_2 & JMP_COND when X"BDB",
            X"BEB" when X"BDC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"BDD",
            X"002" when X"BDE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BDF",
            X"052" when X"BE0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BE1",
            X"051" when X"BE2",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BE3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BE4",
            X"010" when X"BE5",
            X"0" & TYPE_1 & ALU_SUB when X"BE6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BE7",
            X"053" when X"BE8",
            X"0" & TYPE_2 & JMP_UNCOND when X"BE9",
            X"BF7" when X"BEA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"BEB",
            X"001" when X"BEC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BED",
            X"052" when X"BEE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BEF",
            X"051" when X"BF0",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BF1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BF2",
            X"008" when X"BF3",
            X"0" & TYPE_1 & ALU_SUB when X"BF4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BF5",
            X"053" when X"BF6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"BF7",
            X"001" when X"BF8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"BF9",
            X"054" when X"BFA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"BFB",
            X"053" when X"BFC",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"BFD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"BFE",
            X"000" when X"BFF",
            X"0" & TYPE_1 & ALU_CMPE when X"C00",
            X"0" & TYPE_2 & JMP_COND when X"C01",
            X"C16" when X"C02",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C03",
            X"054" when X"C04",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C05",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C06",
            X"000" when X"C07",
            X"0" & TYPE_1 & ALU_ADD when X"C08",
            X"0" & TYPE_1 & ALU_SHIFTL when X"C09",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C0A",
            X"054" when X"C0B",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C0C",
            X"053" when X"C0D",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C0E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C0F",
            X"001" when X"C10",
            X"0" & TYPE_1 & ALU_SUB when X"C11",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C12",
            X"053" when X"C13",
            X"0" & TYPE_2 & JMP_UNCOND when X"C14",
            X"BFB" when X"C15",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C16",
            X"052" when X"C17",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"C18",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"C19",
            X"01B" when X"C1A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C1B",
            X"041" when X"C1C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C1D",
            X"054" when X"C1E",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_B when X"C1F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C20",
            X"041" when X"C21",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C22",
            X"0" & TYPE_1 & ALU_OR when X"C23",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C24",
            X"041" when X"C25",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C26",
            X"052" when X"C27",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"C28",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"C29",
            X"041" when X"C2A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"C2B",
            X"01B" when X"C2C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"C2D",
            X"01A" when X"C2E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C2F",
            X"000" when X"C30",
            X"0" & TYPE_1 & ALU_ADD when X"C31",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C32",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C33",
            X"001" when X"C34",
            X"0" & TYPE_1 & ALU_AND when X"C35",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C36",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C37",
            X"000" when X"C38",
            X"0" & TYPE_1 & ALU_CMPE when X"C39",
            X"0" & TYPE_2 & JMP_COND when X"C3A",
            X"C3E" when X"C3B",
            X"0" & TYPE_2 & JMP_UNCOND when X"C3C",
            X"C42" when X"C3D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C3E",
            X"000" when X"C3F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C40",
            X"049" when X"C41",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"C42",
            X"01A" when X"C43",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C44",
            X"000" when X"C45",
            X"0" & TYPE_1 & ALU_ADD when X"C46",
            X"0" & TYPE_1 & ALU_SHIFTR when X"C47",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C48",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C49",
            X"001" when X"C4A",
            X"0" & TYPE_1 & ALU_AND when X"C4B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"C4C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C4D",
            X"001" when X"C4E",
            X"0" & TYPE_1 & ALU_CMPE when X"C4F",
            X"0" & TYPE_2 & JMP_COND when X"C50",
            X"C54" when X"C51",
            X"0" & TYPE_2 & JMP_UNCOND when X"C52",
            X"DA7" when X"C53",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"C54",
            X"04A" when X"C55",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"C56",
            X"000" when X"C57",
            X"0" & TYPE_1 & ALU_CMPE when X"C58",
            X"0" & TYPE_2 & JMP_COND when X"C59",
            X"C5D" when X"C5A",
            X"0" & TYPE_2 & JMP_UNCOND when X"C5B",
            X"DA7" when X"C5C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C5D",
            X"001" when X"C5E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C5F",
            X"04A" when X"C60",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C61",
            X"042" when X"C62",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C63",
            X"004" when X"C64",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C65",
            X"06F" when X"C66",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C67",
            X"005" when X"C68",
            X"0" & TYPE_4 & I_SEND when X"C69",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C6A",
            X"074" when X"C6B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C6C",
            X"004" when X"C6D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C6E",
            X"06F" when X"C6F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C70",
            X"005" when X"C71",
            X"0" & TYPE_4 & I_SEND when X"C72",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C73",
            X"06E" when X"C74",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C75",
            X"004" when X"C76",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C77",
            X"020" when X"C78",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C79",
            X"005" when X"C7A",
            X"0" & TYPE_4 & I_SEND when X"C7B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C7C",
            X"052" when X"C7D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C7E",
            X"004" when X"C7F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C80",
            X"049" when X"C81",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C82",
            X"005" when X"C83",
            X"0" & TYPE_4 & I_SEND when X"C84",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C85",
            X"047" when X"C86",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C87",
            X"004" when X"C88",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C89",
            X"048" when X"C8A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C8B",
            X"005" when X"C8C",
            X"0" & TYPE_4 & I_SEND when X"C8D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C8E",
            X"054" when X"C8F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C90",
            X"004" when X"C91",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C92",
            X"020" when X"C93",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C94",
            X"005" when X"C95",
            X"0" & TYPE_4 & I_SEND when X"C96",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C97",
            X"070" when X"C98",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C99",
            X"004" when X"C9A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"C9B",
            X"075" when X"C9C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"C9D",
            X"005" when X"C9E",
            X"0" & TYPE_4 & I_SEND when X"C9F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CA0",
            X"06C" when X"CA1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CA2",
            X"004" when X"CA3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CA4",
            X"073" when X"CA5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CA6",
            X"005" when X"CA7",
            X"0" & TYPE_4 & I_SEND when X"CA8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CA9",
            X"061" when X"CAA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CAB",
            X"004" when X"CAC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CAD",
            X"064" when X"CAE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CAF",
            X"005" when X"CB0",
            X"0" & TYPE_4 & I_SEND when X"CB1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CB2",
            X"06F" when X"CB3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CB4",
            X"004" when X"CB5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CB6",
            X"00A" when X"CB7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CB8",
            X"005" when X"CB9",
            X"0" & TYPE_4 & I_SEND when X"CBA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"CBB",
            X"04C" when X"CBC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"CBD",
            X"000" when X"CBE",
            X"0" & TYPE_1 & ALU_CMPG when X"CBF",
            X"0" & TYPE_2 & JMP_COND when X"CC0",
            X"CC4" when X"CC1",
            X"0" & TYPE_2 & JMP_UNCOND when X"CC2",
            X"DA7" when X"CC3",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CC4",
            X"04C" when X"CC5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CC6",
            X"051" when X"CC7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CC8",
            X"000" when X"CC9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CCA",
            X"052" when X"CCB",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CCC",
            X"051" when X"CCD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CCE",
            X"053" when X"CCF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CD0",
            X"051" when X"CD1",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"CD2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"CD3",
            X"008" when X"CD4",
            X"0" & TYPE_1 & ALU_CMPL when X"CD5",
            X"0" & TYPE_2 & JMP_COND when X"CD6",
            X"CFA" when X"CD7",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CD8",
            X"051" when X"CD9",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"CDA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"CDB",
            X"010" when X"CDC",
            X"0" & TYPE_1 & ALU_CMPL when X"CDD",
            X"0" & TYPE_2 & JMP_COND when X"CDE",
            X"CEE" when X"CDF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CE0",
            X"002" when X"CE1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CE2",
            X"052" when X"CE3",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CE4",
            X"051" when X"CE5",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"CE6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"CE7",
            X"010" when X"CE8",
            X"0" & TYPE_1 & ALU_SUB when X"CE9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CEA",
            X"053" when X"CEB",
            X"0" & TYPE_2 & JMP_UNCOND when X"CEC",
            X"CFA" when X"CED",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CEE",
            X"001" when X"CEF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CF0",
            X"052" when X"CF1",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CF2",
            X"051" when X"CF3",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"CF4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"CF5",
            X"008" when X"CF6",
            X"0" & TYPE_1 & ALU_SUB when X"CF7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CF8",
            X"053" when X"CF9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"CFA",
            X"001" when X"CFB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"CFC",
            X"054" when X"CFD",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"CFE",
            X"053" when X"CFF",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D00",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D01",
            X"000" when X"D02",
            X"0" & TYPE_1 & ALU_CMPE when X"D03",
            X"0" & TYPE_2 & JMP_COND when X"D04",
            X"D19" when X"D05",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D06",
            X"054" when X"D07",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D08",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D09",
            X"000" when X"D0A",
            X"0" & TYPE_1 & ALU_ADD when X"D0B",
            X"0" & TYPE_1 & ALU_SHIFTL when X"D0C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D0D",
            X"054" when X"D0E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D0F",
            X"053" when X"D10",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D11",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D12",
            X"001" when X"D13",
            X"0" & TYPE_1 & ALU_SUB when X"D14",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D15",
            X"053" when X"D16",
            X"0" & TYPE_2 & JMP_UNCOND when X"D17",
            X"CFE" when X"D18",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D19",
            X"052" when X"D1A",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"D1B",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"D1C",
            X"01B" when X"D1D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D1E",
            X"041" when X"D1F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D20",
            X"054" when X"D21",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D22",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D23",
            X"0FF" when X"D24",
            X"0" & TYPE_1 & ALU_XOR when X"D25",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_B when X"D26",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D27",
            X"041" when X"D28",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D29",
            X"0" & TYPE_1 & ALU_AND when X"D2A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D2B",
            X"041" when X"D2C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D2D",
            X"052" when X"D2E",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"D2F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D30",
            X"041" when X"D31",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"D32",
            X"01B" when X"D33",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"D34",
            X"04C" when X"D35",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D36",
            X"001" when X"D37",
            X"0" & TYPE_1 & ALU_SUB when X"D38",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D39",
            X"04C" when X"D3A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D3B",
            X"04C" when X"D3C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D3D",
            X"051" when X"D3E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"D3F",
            X"000" when X"D40",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D41",
            X"052" when X"D42",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D43",
            X"051" when X"D44",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D45",
            X"053" when X"D46",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D47",
            X"051" when X"D48",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D49",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D4A",
            X"008" when X"D4B",
            X"0" & TYPE_1 & ALU_CMPL when X"D4C",
            X"0" & TYPE_2 & JMP_COND when X"D4D",
            X"D71" when X"D4E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D4F",
            X"051" when X"D50",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D51",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D52",
            X"010" when X"D53",
            X"0" & TYPE_1 & ALU_CMPL when X"D54",
            X"0" & TYPE_2 & JMP_COND when X"D55",
            X"D65" when X"D56",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"D57",
            X"002" when X"D58",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D59",
            X"052" when X"D5A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D5B",
            X"051" when X"D5C",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D5D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D5E",
            X"010" when X"D5F",
            X"0" & TYPE_1 & ALU_SUB when X"D60",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D61",
            X"053" when X"D62",
            X"0" & TYPE_2 & JMP_UNCOND when X"D63",
            X"D71" when X"D64",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"D65",
            X"001" when X"D66",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D67",
            X"052" when X"D68",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D69",
            X"051" when X"D6A",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D6B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D6C",
            X"008" when X"D6D",
            X"0" & TYPE_1 & ALU_SUB when X"D6E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D6F",
            X"053" when X"D70",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"D71",
            X"001" when X"D72",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D73",
            X"054" when X"D74",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D75",
            X"053" when X"D76",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D77",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D78",
            X"000" when X"D79",
            X"0" & TYPE_1 & ALU_CMPE when X"D7A",
            X"0" & TYPE_2 & JMP_COND when X"D7B",
            X"D90" when X"D7C",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D7D",
            X"054" when X"D7E",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D7F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D80",
            X"000" when X"D81",
            X"0" & TYPE_1 & ALU_ADD when X"D82",
            X"0" & TYPE_1 & ALU_SHIFTL when X"D83",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D84",
            X"054" when X"D85",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D86",
            X"053" when X"D87",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D88",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"D89",
            X"001" when X"D8A",
            X"0" & TYPE_1 & ALU_SUB when X"D8B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D8C",
            X"053" when X"D8D",
            X"0" & TYPE_2 & JMP_UNCOND when X"D8E",
            X"D75" when X"D8F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D90",
            X"052" when X"D91",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"D92",
            X"0" & TYPE_3 & LD & SRC_INDXD_MEM & DST_ACC when X"D93",
            X"01B" when X"D94",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D95",
            X"041" when X"D96",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D97",
            X"054" when X"D98",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_B when X"D99",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"D9A",
            X"041" when X"D9B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"D9C",
            X"0" & TYPE_1 & ALU_OR when X"D9D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"D9E",
            X"041" when X"D9F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"DA0",
            X"052" when X"DA1",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_INDX when X"DA2",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"DA3",
            X"041" when X"DA4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_INDXD_MEM when X"DA5",
            X"01B" when X"DA6",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"DA7",
            X"01A" when X"DA8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DA9",
            X"000" when X"DAA",
            X"0" & TYPE_1 & ALU_ADD when X"DAB",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DAC",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"DAD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DAE",
            X"001" when X"DAF",
            X"0" & TYPE_1 & ALU_AND when X"DB0",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"DB1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DB2",
            X"000" when X"DB3",
            X"0" & TYPE_1 & ALU_CMPE when X"DB4",
            X"0" & TYPE_2 & JMP_COND when X"DB5",
            X"DB9" when X"DB6",
            X"0" & TYPE_2 & JMP_UNCOND when X"DB7",
            X"DBD" when X"DB8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DB9",
            X"000" when X"DBA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DBB",
            X"04A" when X"DBC",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"DBD",
            X"019" when X"DBE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DBF",
            X"000" when X"DC0",
            X"0" & TYPE_1 & ALU_ADD when X"DC1",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC2",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC3",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC4",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC5",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC6",
            X"0" & TYPE_1 & ALU_SHIFTR when X"DC7",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"DC8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DC9",
            X"001" when X"DCA",
            X"0" & TYPE_1 & ALU_AND when X"DCB",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"DCC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DCD",
            X"001" when X"DCE",
            X"0" & TYPE_1 & ALU_CMPE when X"DCF",
            X"0" & TYPE_2 & JMP_COND when X"DD0",
            X"DD4" when X"DD1",
            X"0" & TYPE_2 & JMP_UNCOND when X"DD2",
            X"E85" when X"DD3",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"DD4",
            X"04B" when X"DD5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"DD6",
            X"000" when X"DD7",
            X"0" & TYPE_1 & ALU_CMPE when X"DD8",
            X"0" & TYPE_2 & JMP_COND when X"DD9",
            X"DDD" when X"DDA",
            X"0" & TYPE_2 & JMP_UNCOND when X"DDB",
            X"E85" when X"DDC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DDD",
            X"001" when X"DDE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DDF",
            X"04B" when X"DE0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DE1",
            X"042" when X"DE2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DE3",
            X"004" when X"DE4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DE5",
            X"06F" when X"DE6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DE7",
            X"005" when X"DE8",
            X"0" & TYPE_4 & I_SEND when X"DE9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DEA",
            X"074" when X"DEB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DEC",
            X"004" when X"DED",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DEE",
            X"06F" when X"DEF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DF0",
            X"005" when X"DF1",
            X"0" & TYPE_4 & I_SEND when X"DF2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DF3",
            X"06E" when X"DF4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DF5",
            X"004" when X"DF6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DF7",
            X"020" when X"DF8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DF9",
            X"005" when X"DFA",
            X"0" & TYPE_4 & I_SEND when X"DFB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"DFC",
            X"043" when X"DFD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"DFE",
            X"004" when X"DFF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E00",
            X"045" when X"E01",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E02",
            X"005" when X"E03",
            X"0" & TYPE_4 & I_SEND when X"E04",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E05",
            X"04E" when X"E06",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E07",
            X"004" when X"E08",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E09",
            X"054" when X"E0A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E0B",
            X"005" when X"E0C",
            X"0" & TYPE_4 & I_SEND when X"E0D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E0E",
            X"045" when X"E0F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E10",
            X"004" when X"E11",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E12",
            X"052" when X"E13",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E14",
            X"005" when X"E15",
            X"0" & TYPE_4 & I_SEND when X"E16",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E17",
            X"020" when X"E18",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E19",
            X"004" when X"E1A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E1B",
            X"070" when X"E1C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E1D",
            X"005" when X"E1E",
            X"0" & TYPE_4 & I_SEND when X"E1F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E20",
            X"075" when X"E21",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E22",
            X"004" when X"E23",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E24",
            X"06C" when X"E25",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E26",
            X"005" when X"E27",
            X"0" & TYPE_4 & I_SEND when X"E28",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E29",
            X"073" when X"E2A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E2B",
            X"004" when X"E2C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E2D",
            X"061" when X"E2E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E2F",
            X"005" when X"E30",
            X"0" & TYPE_4 & I_SEND when X"E31",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E32",
            X"064" when X"E33",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E34",
            X"004" when X"E35",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E36",
            X"06F" when X"E37",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E38",
            X"005" when X"E39",
            X"0" & TYPE_4 & I_SEND when X"E3A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E3B",
            X"00A" when X"E3C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E3D",
            X"004" when X"E3E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E3F",
            X"020" when X"E40",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E41",
            X"005" when X"E42",
            X"0" & TYPE_4 & I_SEND when X"E43",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E44",
            X"06C" when X"E45",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E46",
            X"004" when X"E47",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E48",
            X"065" when X"E49",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E4A",
            X"005" when X"E4B",
            X"0" & TYPE_4 & I_SEND when X"E4C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E4D",
            X"064" when X"E4E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E4F",
            X"004" when X"E50",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E51",
            X"05F" when X"E52",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E53",
            X"005" when X"E54",
            X"0" & TYPE_4 & I_SEND when X"E55",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E56",
            X"073" when X"E57",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E58",
            X"004" when X"E59",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E5A",
            X"074" when X"E5B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E5C",
            X"005" when X"E5D",
            X"0" & TYPE_4 & I_SEND when X"E5E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E5F",
            X"061" when X"E60",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E61",
            X"004" when X"E62",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E63",
            X"074" when X"E64",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E65",
            X"005" when X"E66",
            X"0" & TYPE_4 & I_SEND when X"E67",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E68",
            X"065" when X"E69",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E6A",
            X"004" when X"E6B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E6C",
            X"03A" when X"E6D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E6E",
            X"005" when X"E6F",
            X"0" & TYPE_4 & I_SEND when X"E70",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E71",
            X"020" when X"E72",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E73",
            X"004" when X"E74",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"E75",
            X"04C" when X"E76",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"E77",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"E78",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E79",
            X"005" when X"E7A",
            X"0" & TYPE_4 & I_SEND when X"E7B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E7C",
            X"00A" when X"E7D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E7E",
            X"004" when X"E7F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E80",
            X"020" when X"E81",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E82",
            X"005" when X"E83",
            X"0" & TYPE_4 & I_SEND when X"E84",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"E85",
            X"019" when X"E86",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"E87",
            X"000" when X"E88",
            X"0" & TYPE_1 & ALU_ADD when X"E89",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8A",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8B",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8C",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8D",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8E",
            X"0" & TYPE_1 & ALU_SHIFTR when X"E8F",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"E90",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"E91",
            X"001" when X"E92",
            X"0" & TYPE_1 & ALU_AND when X"E93",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"E94",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"E95",
            X"000" when X"E96",
            X"0" & TYPE_1 & ALU_CMPE when X"E97",
            X"0" & TYPE_2 & JMP_COND when X"E98",
            X"E9C" when X"E99",
            X"0" & TYPE_2 & JMP_UNCOND when X"E9A",
            X"EA0" when X"E9B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"E9C",
            X"000" when X"E9D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"E9E",
            X"04B" when X"E9F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EA0",
            X"018" when X"EA1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EA2",
            X"000" when X"EA3",
            X"0" & TYPE_1 & ALU_ADD when X"EA4",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EA5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EA6",
            X"001" when X"EA7",
            X"0" & TYPE_1 & ALU_AND when X"EA8",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EA9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EAA",
            X"000" when X"EAB",
            X"0" & TYPE_1 & ALU_CMPE when X"EAC",
            X"0" & TYPE_2 & JMP_COND when X"EAD",
            X"EB8" when X"EAE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EAF",
            X"01C" when X"EB0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EB1",
            X"001" when X"EB2",
            X"0" & TYPE_1 & ALU_OR when X"EB3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"EB4",
            X"01C" when X"EB5",
            X"0" & TYPE_2 & JMP_UNCOND when X"EB6",
            X"EBF" when X"EB7",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EB8",
            X"01C" when X"EB9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EBA",
            X"0FE" when X"EBB",
            X"0" & TYPE_1 & ALU_AND when X"EBC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"EBD",
            X"01C" when X"EBE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EBF",
            X"018" when X"EC0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EC1",
            X"000" when X"EC2",
            X"0" & TYPE_1 & ALU_ADD when X"EC3",
            X"0" & TYPE_1 & ALU_SHIFTR when X"EC4",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EC5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EC6",
            X"001" when X"EC7",
            X"0" & TYPE_1 & ALU_AND when X"EC8",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EC9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ECA",
            X"000" when X"ECB",
            X"0" & TYPE_1 & ALU_CMPE when X"ECC",
            X"0" & TYPE_2 & JMP_COND when X"ECD",
            X"ED8" when X"ECE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"ECF",
            X"01C" when X"ED0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"ED1",
            X"002" when X"ED2",
            X"0" & TYPE_1 & ALU_OR when X"ED3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"ED4",
            X"01C" when X"ED5",
            X"0" & TYPE_2 & JMP_UNCOND when X"ED6",
            X"EDF" when X"ED7",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"ED8",
            X"01C" when X"ED9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EDA",
            X"0FD" when X"EDB",
            X"0" & TYPE_1 & ALU_AND when X"EDC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"EDD",
            X"01C" when X"EDE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EDF",
            X"018" when X"EE0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EE1",
            X"000" when X"EE2",
            X"0" & TYPE_1 & ALU_ADD when X"EE3",
            X"0" & TYPE_1 & ALU_SHIFTR when X"EE4",
            X"0" & TYPE_1 & ALU_SHIFTR when X"EE5",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EE6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EE7",
            X"001" when X"EE8",
            X"0" & TYPE_1 & ALU_AND when X"EE9",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"EEA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EEB",
            X"000" when X"EEC",
            X"0" & TYPE_1 & ALU_CMPE when X"EED",
            X"0" & TYPE_2 & JMP_COND when X"EEE",
            X"EF9" when X"EEF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EF0",
            X"01C" when X"EF1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EF2",
            X"004" when X"EF3",
            X"0" & TYPE_1 & ALU_OR when X"EF4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"EF5",
            X"01C" when X"EF6",
            X"0" & TYPE_2 & JMP_UNCOND when X"EF7",
            X"F00" when X"EF8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"EF9",
            X"01C" when X"EFA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"EFB",
            X"0FB" when X"EFC",
            X"0" & TYPE_1 & ALU_AND when X"EFD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"EFE",
            X"01C" when X"EFF",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F00",
            X"018" when X"F01",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F02",
            X"000" when X"F03",
            X"0" & TYPE_1 & ALU_ADD when X"F04",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F05",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F06",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F07",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F08",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F09",
            X"001" when X"F0A",
            X"0" & TYPE_1 & ALU_AND when X"F0B",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F0C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F0D",
            X"000" when X"F0E",
            X"0" & TYPE_1 & ALU_CMPE when X"F0F",
            X"0" & TYPE_2 & JMP_COND when X"F10",
            X"F1B" when X"F11",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F12",
            X"01C" when X"F13",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F14",
            X"008" when X"F15",
            X"0" & TYPE_1 & ALU_OR when X"F16",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F17",
            X"01C" when X"F18",
            X"0" & TYPE_2 & JMP_UNCOND when X"F19",
            X"F22" when X"F1A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F1B",
            X"01C" when X"F1C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F1D",
            X"0F7" when X"F1E",
            X"0" & TYPE_1 & ALU_AND when X"F1F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F20",
            X"01C" when X"F21",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F22",
            X"018" when X"F23",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F24",
            X"000" when X"F25",
            X"0" & TYPE_1 & ALU_ADD when X"F26",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F27",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F28",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F29",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F2A",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F2B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F2C",
            X"001" when X"F2D",
            X"0" & TYPE_1 & ALU_AND when X"F2E",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F2F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F30",
            X"000" when X"F31",
            X"0" & TYPE_1 & ALU_CMPE when X"F32",
            X"0" & TYPE_2 & JMP_COND when X"F33",
            X"F3E" when X"F34",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F35",
            X"01C" when X"F36",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F37",
            X"010" when X"F38",
            X"0" & TYPE_1 & ALU_OR when X"F39",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F3A",
            X"01C" when X"F3B",
            X"0" & TYPE_2 & JMP_UNCOND when X"F3C",
            X"F45" when X"F3D",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F3E",
            X"01C" when X"F3F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F40",
            X"0EF" when X"F41",
            X"0" & TYPE_1 & ALU_AND when X"F42",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F43",
            X"01C" when X"F44",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F45",
            X"018" when X"F46",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F47",
            X"000" when X"F48",
            X"0" & TYPE_1 & ALU_ADD when X"F49",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F4A",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F4B",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F4C",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F4D",
            X"0" & TYPE_1 & ALU_SHIFTR when X"F4E",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F4F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F50",
            X"001" when X"F51",
            X"0" & TYPE_1 & ALU_AND when X"F52",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"F53",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F54",
            X"000" when X"F55",
            X"0" & TYPE_1 & ALU_CMPE when X"F56",
            X"0" & TYPE_2 & JMP_COND when X"F57",
            X"F62" when X"F58",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F59",
            X"01C" when X"F5A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F5B",
            X"020" when X"F5C",
            X"0" & TYPE_1 & ALU_OR when X"F5D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F5E",
            X"01C" when X"F5F",
            X"0" & TYPE_2 & JMP_UNCOND when X"F60",
            X"F69" when X"F61",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"F62",
            X"01C" when X"F63",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"F64",
            X"0DF" when X"F65",
            X"0" & TYPE_1 & ALU_AND when X"F66",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"F67",
            X"01C" when X"F68",
            X"0" & TYPE_2 & JMP_UNCOND when X"F69",
            X"958" when X"F6A",
            X"0" & TYPE_1 & ALU_ADD when others;
end AUTOMATIC;