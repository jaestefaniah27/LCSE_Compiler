LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE work.PIC_pkg.all;

entity ROM_Generated is
  port (
    Instruction     : out std_logic_vector(11 downto 0);
    Program_counter : in  std_logic_vector(11 downto 0));
end ROM_Generated;

architecture AUTOMATIC of ROM_Generated is
begin
    with Program_counter select
        Instruction <=
            X"0" & TYPE_2 & JMP_UNCOND when X"000",
            X"003" when X"001",
            X"0" & TYPE_4 & I_RETI when X"002",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"003",
            X"000" when X"004",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"005",
            X"050" when X"006",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"007",
            X"001" when X"008",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"009",
            X"051" when X"00A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"00B",
            X"000" when X"00C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"00D",
            X"052" when X"00E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"00F",
            X"000" when X"010",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"011",
            X"053" when X"012",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"013",
            X"001" when X"014",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"015",
            X"05B" when X"016",
            X"0" & TYPE_2 & JMP_UNCOND when X"017",
            X"019" when X"018",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"019",
            X"053" when X"01A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"01B",
            X"004" when X"01C",
            X"0" & TYPE_4 & I_SEND when X"01D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"01E",
            X"049" when X"01F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"020",
            X"004" when X"021",
            X"0" & TYPE_4 & I_SEND when X"022",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"023",
            X"053" when X"024",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"025",
            X"004" when X"026",
            X"0" & TYPE_4 & I_SEND when X"027",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"028",
            X"054" when X"029",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"02A",
            X"004" when X"02B",
            X"0" & TYPE_4 & I_SEND when X"02C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"02D",
            X"045" when X"02E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"02F",
            X"004" when X"030",
            X"0" & TYPE_4 & I_SEND when X"031",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"032",
            X"04D" when X"033",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"034",
            X"004" when X"035",
            X"0" & TYPE_4 & I_SEND when X"036",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"037",
            X"041" when X"038",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"039",
            X"004" when X"03A",
            X"0" & TYPE_4 & I_SEND when X"03B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"03C",
            X"020" when X"03D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"03E",
            X"004" when X"03F",
            X"0" & TYPE_4 & I_SEND when X"040",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"041",
            X"04C" when X"042",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"043",
            X"004" when X"044",
            X"0" & TYPE_4 & I_SEND when X"045",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"046",
            X"049" when X"047",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"048",
            X"004" when X"049",
            X"0" & TYPE_4 & I_SEND when X"04A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"04B",
            X"053" when X"04C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"04D",
            X"004" when X"04E",
            X"0" & TYPE_4 & I_SEND when X"04F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"050",
            X"054" when X"051",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"052",
            X"004" when X"053",
            X"0" & TYPE_4 & I_SEND when X"054",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"055",
            X"04F" when X"056",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"057",
            X"004" when X"058",
            X"0" & TYPE_4 & I_SEND when X"059",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"05A",
            X"03A" when X"05B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"05C",
            X"004" when X"05D",
            X"0" & TYPE_4 & I_SEND when X"05E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"05F",
            X"020" when X"060",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"061",
            X"004" when X"062",
            X"0" & TYPE_4 & I_SEND when X"063",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"064",
            X"046" when X"065",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"066",
            X"004" when X"067",
            X"0" & TYPE_4 & I_SEND when X"068",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"069",
            X"049" when X"06A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"06B",
            X"004" when X"06C",
            X"0" & TYPE_4 & I_SEND when X"06D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"06E",
            X"042" when X"06F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"070",
            X"004" when X"071",
            X"0" & TYPE_4 & I_SEND when X"072",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"073",
            X"04F" when X"074",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"075",
            X"004" when X"076",
            X"0" & TYPE_4 & I_SEND when X"077",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"078",
            X"04E" when X"079",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"07A",
            X"004" when X"07B",
            X"0" & TYPE_4 & I_SEND when X"07C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"07D",
            X"041" when X"07E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"07F",
            X"004" when X"080",
            X"0" & TYPE_4 & I_SEND when X"081",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"082",
            X"043" when X"083",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"084",
            X"004" when X"085",
            X"0" & TYPE_4 & I_SEND when X"086",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"087",
            X"043" when X"088",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"089",
            X"004" when X"08A",
            X"0" & TYPE_4 & I_SEND when X"08B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"08C",
            X"049" when X"08D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"08E",
            X"004" when X"08F",
            X"0" & TYPE_4 & I_SEND when X"090",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"091",
            X"020" when X"092",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"093",
            X"004" when X"094",
            X"0" & TYPE_4 & I_SEND when X"095",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"096",
            X"028" when X"097",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"098",
            X"004" when X"099",
            X"0" & TYPE_4 & I_SEND when X"09A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"09B",
            X"046" when X"09C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"09D",
            X"004" when X"09E",
            X"0" & TYPE_4 & I_SEND when X"09F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0A0",
            X"06C" when X"0A1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0A2",
            X"004" when X"0A3",
            X"0" & TYPE_4 & I_SEND when X"0A4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0A5",
            X"061" when X"0A6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0A7",
            X"004" when X"0A8",
            X"0" & TYPE_4 & I_SEND when X"0A9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0AA",
            X"06E" when X"0AB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0AC",
            X"004" when X"0AD",
            X"0" & TYPE_4 & I_SEND when X"0AE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0AF",
            X"063" when X"0B0",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0B1",
            X"004" when X"0B2",
            X"0" & TYPE_4 & I_SEND when X"0B3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0B4",
            X"06F" when X"0B5",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0B6",
            X"004" when X"0B7",
            X"0" & TYPE_4 & I_SEND when X"0B8",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0B9",
            X"073" when X"0BA",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0BB",
            X"004" when X"0BC",
            X"0" & TYPE_4 & I_SEND when X"0BD",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0BE",
            X"029" when X"0BF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0C0",
            X"004" when X"0C1",
            X"0" & TYPE_4 & I_SEND when X"0C2",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0C3",
            X"02E" when X"0C4",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0C5",
            X"004" when X"0C6",
            X"0" & TYPE_4 & I_SEND when X"0C7",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0C8",
            X"020" when X"0C9",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0CA",
            X"004" when X"0CB",
            X"0" & TYPE_4 & I_SEND when X"0CC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0CD",
            X"050" when X"0CE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0CF",
            X"004" when X"0D0",
            X"0" & TYPE_4 & I_SEND when X"0D1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0D2",
            X"055" when X"0D3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0D4",
            X"004" when X"0D5",
            X"0" & TYPE_4 & I_SEND when X"0D6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0D7",
            X"04C" when X"0D8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0D9",
            X"004" when X"0DA",
            X"0" & TYPE_4 & I_SEND when X"0DB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0DC",
            X"053" when X"0DD",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0DE",
            X"004" when X"0DF",
            X"0" & TYPE_4 & I_SEND when X"0E0",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0E1",
            X"041" when X"0E2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0E3",
            X"004" when X"0E4",
            X"0" & TYPE_4 & I_SEND when X"0E5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0E6",
            X"052" when X"0E7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0E8",
            X"004" when X"0E9",
            X"0" & TYPE_4 & I_SEND when X"0EA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0EB",
            X"020" when X"0EC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0ED",
            X"004" when X"0EE",
            X"0" & TYPE_4 & I_SEND when X"0EF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0F0",
            X"043" when X"0F1",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0F2",
            X"004" when X"0F3",
            X"0" & TYPE_4 & I_SEND when X"0F4",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0F5",
            X"045" when X"0F6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0F7",
            X"004" when X"0F8",
            X"0" & TYPE_4 & I_SEND when X"0F9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0FA",
            X"04E" when X"0FB",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"0FC",
            X"004" when X"0FD",
            X"0" & TYPE_4 & I_SEND when X"0FE",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"0FF",
            X"054" when X"100",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"101",
            X"004" when X"102",
            X"0" & TYPE_4 & I_SEND when X"103",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"104",
            X"052" when X"105",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"106",
            X"004" when X"107",
            X"0" & TYPE_4 & I_SEND when X"108",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"109",
            X"041" when X"10A",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"10B",
            X"004" when X"10C",
            X"0" & TYPE_4 & I_SEND when X"10D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"10E",
            X"04C" when X"10F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"110",
            X"004" when X"111",
            X"0" & TYPE_4 & I_SEND when X"112",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"113",
            X"00A" when X"114",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"115",
            X"004" when X"116",
            X"0" & TYPE_4 & I_SEND when X"117",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"118",
            X"054" when X"119",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"11A",
            X"055" when X"11B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"11C",
            X"001" when X"11D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"11E",
            X"056" when X"11F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"120",
            X"055" when X"121",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"122",
            X"056" when X"123",
            X"0" & TYPE_1 & ALU_CMPE when X"124",
            X"0" & TYPE_2 & JMP_COND when X"125",
            X"12B" when X"126",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"127",
            X"000" when X"128",
            X"0" & TYPE_2 & JMP_UNCOND when X"129",
            X"12D" when X"12A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"12B",
            X"001" when X"12C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"12D",
            X"057" when X"12E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"12F",
            X"053" when X"130",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"131",
            X"058" when X"132",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"133",
            X"000" when X"134",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"135",
            X"059" when X"136",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"137",
            X"058" when X"138",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"139",
            X"059" when X"13A",
            X"0" & TYPE_1 & ALU_CMPE when X"13B",
            X"0" & TYPE_2 & JMP_COND when X"13C",
            X"142" when X"13D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"13E",
            X"000" when X"13F",
            X"0" & TYPE_2 & JMP_UNCOND when X"140",
            X"144" when X"141",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"142",
            X"001" when X"143",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"144",
            X"05A" when X"145",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"146",
            X"057" when X"147",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"148",
            X"05A" when X"149",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"14A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"14B",
            X"000" when X"14C",
            X"0" & TYPE_1 & ALU_CMPE when X"14D",
            X"0" & TYPE_2 & JMP_COND when X"14E",
            X"235" when X"14F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"150",
            X"000" when X"151",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"152",
            X"050" when X"153",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"154",
            X"001" when X"155",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"156",
            X"051" when X"157",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"158",
            X"053" when X"159",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"15A",
            X"004" when X"15B",
            X"0" & TYPE_4 & I_SEND when X"15C",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"15D",
            X"065" when X"15E",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"15F",
            X"004" when X"160",
            X"0" & TYPE_4 & I_SEND when X"161",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"162",
            X"063" when X"163",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"164",
            X"004" when X"165",
            X"0" & TYPE_4 & I_SEND when X"166",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"167",
            X"075" when X"168",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"169",
            X"004" when X"16A",
            X"0" & TYPE_4 & I_SEND when X"16B",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"16C",
            X"065" when X"16D",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"16E",
            X"004" when X"16F",
            X"0" & TYPE_4 & I_SEND when X"170",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"171",
            X"06E" when X"172",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"173",
            X"004" when X"174",
            X"0" & TYPE_4 & I_SEND when X"175",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"176",
            X"063" when X"177",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"178",
            X"004" when X"179",
            X"0" & TYPE_4 & I_SEND when X"17A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"17B",
            X"069" when X"17C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"17D",
            X"004" when X"17E",
            X"0" & TYPE_4 & I_SEND when X"17F",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"180",
            X"061" when X"181",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"182",
            X"004" when X"183",
            X"0" & TYPE_4 & I_SEND when X"184",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"185",
            X"03A" when X"186",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"187",
            X"004" when X"188",
            X"0" & TYPE_4 & I_SEND when X"189",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"18A",
            X"020" when X"18B",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"18C",
            X"004" when X"18D",
            X"0" & TYPE_4 & I_SEND when X"18E",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"18F",
            X"050" when X"190",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"191",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"192",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"193",
            X"004" when X"194",
            X"0" & TYPE_4 & I_SEND when X"195",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"196",
            X"02C" when X"197",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"198",
            X"004" when X"199",
            X"0" & TYPE_4 & I_SEND when X"19A",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"19B",
            X"020" when X"19C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"19D",
            X"004" when X"19E",
            X"0" & TYPE_4 & I_SEND when X"19F",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1A0",
            X"051" when X"1A1",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"1A2",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"1A3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1A4",
            X"004" when X"1A5",
            X"0" & TYPE_4 & I_SEND when X"1A6",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1A7",
            X"05B" when X"1A8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1A9",
            X"05C" when X"1AA",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1AB",
            X"001" when X"1AC",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1AD",
            X"05D" when X"1AE",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1AF",
            X"05C" when X"1B0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"1B1",
            X"05D" when X"1B2",
            X"0" & TYPE_1 & ALU_CMPE when X"1B3",
            X"0" & TYPE_2 & JMP_COND when X"1B4",
            X"1BA" when X"1B5",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1B6",
            X"000" when X"1B7",
            X"0" & TYPE_2 & JMP_UNCOND when X"1B8",
            X"1BC" when X"1B9",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1BA",
            X"001" when X"1BB",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"1BC",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"1BD",
            X"000" when X"1BE",
            X"0" & TYPE_1 & ALU_CMPE when X"1BF",
            X"0" & TYPE_2 & JMP_COND when X"1C0",
            X"22E" when X"1C1",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1C2",
            X"050" when X"1C3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1C4",
            X"05E" when X"1C5",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1C6",
            X"051" when X"1C7",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1C8",
            X"05F" when X"1C9",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1CA",
            X"05E" when X"1CB",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"1CC",
            X"05F" when X"1CD",
            X"0" & TYPE_1 & ALU_ADD when X"1CE",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1CF",
            X"052" when X"1D0",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1D1",
            X"052" when X"1D2",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1D3",
            X"060" when X"1D4",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1D5",
            X"050" when X"1D6",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1D7",
            X"061" when X"1D8",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"1D9",
            X"060" when X"1DA",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"1DB",
            X"061" when X"1DC",
            X"0" & TYPE_1 & ALU_CMPL when X"1DD",
            X"0" & TYPE_2 & JMP_COND when X"1DE",
            X"1E4" when X"1DF",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1E0",
            X"000" when X"1E1",
            X"0" & TYPE_2 & JMP_UNCOND when X"1E2",
            X"1E6" when X"1E3",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1E4",
            X"001" when X"1E5",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"1E6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"1E7",
            X"000" when X"1E8",
            X"0" & TYPE_1 & ALU_CMPE when X"1E9",
            X"0" & TYPE_2 & JMP_COND when X"1EA",
            X"1F2" when X"1EB",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1EC",
            X"000" when X"1ED",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1EE",
            X"05B" when X"1EF",
            X"0" & TYPE_2 & JMP_UNCOND when X"1F0",
            X"22C" when X"1F1",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1F2",
            X"02C" when X"1F3",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1F4",
            X"004" when X"1F5",
            X"0" & TYPE_4 & I_SEND when X"1F6",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"1F7",
            X"020" when X"1F8",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"1F9",
            X"004" when X"1FA",
            X"0" & TYPE_4 & I_SEND when X"1FB",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"1FC",
            X"052" when X"1FD",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"1FE",
            X"0" & TYPE_1 & ALU_BIN2ASCII when X"1FF",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"200",
            X"004" when X"201",
            X"0" & TYPE_4 & I_SEND when X"202",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"203",
            X"051" when X"204",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"205",
            X"050" when X"206",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"207",
            X"052" when X"208",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"209",
            X"051" when X"20A",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"20B",
            X"050" when X"20C",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"20D",
            X"062" when X"20E",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"20F",
            X"090" when X"210",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"211",
            X"063" when X"212",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_A when X"213",
            X"062" when X"214",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_B when X"215",
            X"063" when X"216",
            X"0" & TYPE_1 & ALU_CMPG when X"217",
            X"0" & TYPE_2 & JMP_COND when X"218",
            X"21E" when X"219",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"21A",
            X"000" when X"21B",
            X"0" & TYPE_2 & JMP_UNCOND when X"21C",
            X"220" when X"21D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"21E",
            X"001" when X"21F",
            X"0" & TYPE_3 & LD & SRC_ACC & DST_A when X"220",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_B when X"221",
            X"000" when X"222",
            X"0" & TYPE_1 & ALU_CMPE when X"223",
            X"0" & TYPE_2 & JMP_COND when X"224",
            X"22C" when X"225",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"226",
            X"000" when X"227",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"228",
            X"05B" when X"229",
            X"0" & TYPE_2 & JMP_UNCOND when X"22A",
            X"22C" when X"22B",
            X"0" & TYPE_2 & JMP_UNCOND when X"22C",
            X"1A7" when X"22D",
            X"0" & TYPE_3 & LD & SRC_CONSTANT & DST_ACC when X"22E",
            X"00A" when X"22F",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"230",
            X"004" when X"231",
            X"0" & TYPE_4 & I_SEND when X"232",
            X"0" & TYPE_2 & JMP_UNCOND when X"233",
            X"235" when X"234",
            X"0" & TYPE_3 & LD & SRC_MEM & DST_ACC when X"235",
            X"054" when X"236",
            X"0" & TYPE_3 & WR & SRC_ACC & DST_MEM when X"237",
            X"053" when X"238",
            X"0" & TYPE_2 & JMP_UNCOND when X"239",
            X"118" when X"23A",
            X"0" & TYPE_1 & ALU_ADD when others;
end AUTOMATIC;